netcdf ATL08_20181014084920_02400109_003_01 {
dimensions:
	ds_geosegments = 5 ;
	ds_metrics = 9 ;
	ds_surf_type = 5 ;
variables:
	byte ds_geosegments(ds_geosegments) ;
		ds_geosegments:long_name = "Geosegments" ;
		ds_geosegments:units = "1" ;
		ds_geosegments:valid_min = 1b ;
		ds_geosegments:valid_max = 5b ;
		ds_geosegments:flag_values = 1b, 2b, 3b, 4b, 5b ;
		ds_geosegments:flag_meanings = "geosegments1 geosegments2 geosegments3 geosegments4 geosegments5" ;
		ds_geosegments:description = "Dimension scale for geosegments within land segments." ;
	byte ds_metrics(ds_metrics) ;
		ds_metrics:contentType = "referenceInformation" ;
		ds_metrics:description = "Dimension scale for metrics." ;
		ds_metrics:flag_meanings = "metrics1 metrics2 metrics3 metrics4 metrics5 metrics6 metrics7 metrics8 metrics9" ;
		ds_metrics:flag_values = 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		ds_metrics:long_name = "Metrics" ;
		ds_metrics:units = "1" ;
		ds_metrics:valid_max = 4b ;
		ds_metrics:valid_min = 1b ;
	int ds_surf_type(ds_surf_type) ;
		ds_surf_type:contentType = "auxiliaryInformation" ;
		ds_surf_type:units = "1" ;
		ds_surf_type:description = "Dimension scale indexing the surface type array. Index=1 corresponds to Land; index = 2 corresponds to Ocean; Index = 3 corresponds to SeaIce; Index=4 corresponds to LandIce; Index=5 corresponds to InlandWater" ;
		ds_surf_type:flag_meanings = "land ocean seaice landice inland_water" ;
		ds_surf_type:flag_values = 1, 2, 3, 4, 5 ;
		ds_surf_type:long_name = "Surface Type Dimension Scale" ;
		ds_surf_type:valid_max = 5 ;
		ds_surf_type:valid_min = 1 ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:contributor_name = "Thomas E Neumann (thomas.neumann@nasa.gov), Thorsten Markus (thorsten.markus@nasa.gov), Suneel Bhardwaj (suneel.bhardwaj@nasa.gov) David W Hancock III (david.w.hancock@nasa.gov)" ;
		:contributor_role = "Instrument Engineer, Investigator, Principle Investigator, Data Producer, Data Producer" ;
		:date_type = "UTC" ;
		:description = "This data set (ATL08) contains along-track heights above the WGS84 ellipsoid (ITRF2014 reference frame) for the ground and canopy surfaces. The canopy and ground surfaces are processed in fixed 100 m data segments, which typically contain more than 100 sig" ;
		:featureType = "trajectory" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:granule_type = "ATL08" ;
		:identifier_product_doi_authority = "http://dx.doi.org" ;
		:level = "L3A" ;
		:license = "Data may not be reproduced or distributed without including the citation for this product included in this metadata. Data may not be distributed in an altered form without the written permission of the ICESat-2 Science Project Office at NASA/GSFC." ;
		:naming_authority = "http://dx.doi.org" ;
		:short_name = "ATL08" ;
		:spatial_coverage_type = "Horizontal" ;
		:standard_name_vocabulary = "CF-1.6" ;
		:time_type = "CCSDS UTC-A" ;
		:title = "SET_BY_META" ;
		:date_created = "2020-04-01T14:03:26.000000Z" ;
		:hdfversion = "HDF5 1.10.3" ;
		:history = "2020-04-01T14:03:26.000000Z;ae899cbd-cf20-3541-9952-cb5220d5467b;Created by PGE atlas_l3a_ld Version 3.3.1" ;
		:identifier_file_uuid = "ae899cbd-cf20-3541-9952-cb5220d5467b" ;
		:identifier_product_format_version = "3.3" ;
		:time_coverage_duration = 362. ;
		:time_coverage_end = "2018-10-14T08:55:22.000000Z" ;
		:time_coverage_start = "2018-10-14T08:49:20.000000Z" ;
		:geospatial_lat_min = -33.6709309916173 ;
		:geospatial_lon_min = -80.4279359434023 ;
		:geospatial_lat_max = -33.6666200966049 ;
		:geospatial_lon_max = -80.4274386927379 ;
		:publisher_name = "NSIDC DAAC > NASA National Snow and Ice Data Center Distributed Active Archive Center" ;
		:publisher_email = "nsidc@nsidc.org" ;
		:publisher_url = "http://nsidc.org/daac/" ;
		:identifier_product_type = "ATL08" ;
		:identifier_product_doi = "doi:10.5067/ATLAS/ATL08.003" ;
		:institution = "National Aeronautics and Space Administration (NASA)" ;
		:creator_name = "GSFC I-SIPS > ICESat-2 Science Investigator-led Processing System" ;
		:summary = "The purpose of ATL08 is to provide along-track land/canopy heights and associated statistics." ;
		:keywords = "EARTH SCIENCE > BIOSPHERE > VEGETATION > NONE > NONE > NONE > NONE" ;
		:keywords_vocabulary = "NASA/GCMD Science Keywords" ;
		:citation = "Cite these data in publications as follows: The data used in this study were produced by the ICESat-2 Science Project Office at NASA/GSFC. The data archive site is the NASA National Snow and Ice Data Center Distributed Active Archive Center." ;
		:processing_level = "3A" ;
		:references = "http://nsidc.org/data/icesat2/data.html" ;
		:project = "ICESat-2 > Ice, Cloud, and land Elevation Satellite-2" ;
		:instrument = "ATLAS > Advanced Topographic Laser Altimeter System" ;
		:platform = "ICESat-2 > Ice, Cloud, and land Elevation Satellite-2" ;
		:source = "Spacecraft" ;

group: ancillary_data {
  dimensions:
  	phony_dim_9 = 1 ;
  variables:
  	double atlas_sdp_gps_epoch(phony_dim_9) ;
  		atlas_sdp_gps_epoch:contentType = "auxiliaryInformation" ;
  		atlas_sdp_gps_epoch:description = "Number of GPS seconds between the GPS epoch (1980-01-06T00:00:00.000000Z UTC) and the ATLAS Standard Data Product (SDP) epoch (2018-01-01:T00.00.00.000000 UTC). Add this value to delta time parameters to compute full gps_seconds (relative to the GPS epoch) for each data point." ;
  		atlas_sdp_gps_epoch:long_name = "ATLAS Epoch Offset" ;
  		atlas_sdp_gps_epoch:source = "Operations" ;
  		atlas_sdp_gps_epoch:units = "seconds since 1980-01-06T00:00:00.000000Z" ;
  	string control(phony_dim_9) ;
  		control:contentType = "auxiliaryInformation" ;
  		control:description = "PGE-specific control file used to generate this granule. To re-use, replace breaks (BR) with linefeeds." ;
  		control:long_name = "Control File" ;
  		control:source = "Operations" ;
  		control:units = "1" ;
  	string data_end_utc(phony_dim_9) ;
  		data_end_utc:contentType = "auxiliaryInformation" ;
  		data_end_utc:description = "UTC (in CCSDS-A format) of the last data point within the granule." ;
  		data_end_utc:long_name = "End UTC Time of Granule (CCSDS-A, Actual)" ;
  		data_end_utc:source = "Derived" ;
  		data_end_utc:units = "1" ;
  	string data_start_utc(phony_dim_9) ;
  		data_start_utc:contentType = "auxiliaryInformation" ;
  		data_start_utc:description = "UTC (in CCSDS-A format) of the first data point within the granule." ;
  		data_start_utc:long_name = "Start UTC Time of Granule (CCSDS-A, Actual)" ;
  		data_start_utc:source = "Derived" ;
  		data_start_utc:units = "1" ;
  	int end_cycle(phony_dim_9) ;
  		end_cycle:contentType = "auxiliaryInformation" ;
  		end_cycle:description = "The ending cycle number associated with the data contained within this granule. The cycle number is the counter of the number of 91-day repeat cycles completed by the mission." ;
  		end_cycle:long_name = "Ending Cycle" ;
  		end_cycle:source = "Derived" ;
  		end_cycle:units = "1" ;
  		end_cycle:valid_max = 99 ;
  		end_cycle:valid_min = 0 ;
  	double end_delta_time(phony_dim_9) ;
  		end_delta_time:contentType = "auxiliaryInformation" ;
  		end_delta_time:description = "Number of GPS seconds since the ATLAS SDP epoch at the last data point in the file. The ATLAS Standard Data Products (SDP) epoch offset is defined within /ancillary_data/atlas_sdp_gps_epoch as the number of GPS seconds between the GPS epoch (1980-01-06T00:00:00.000000Z UTC) and the ATLAS SDP epoch. By adding the offset contained within atlas_sdp_gps_epoch to delta time parameters, the time in gps_seconds relative to the GPS epoch can be computed." ;
  		end_delta_time:long_name = "ATLAS End Time (Actual)" ;
  		end_delta_time:source = "Derived" ;
  		end_delta_time:standard_name = "time" ;
  		end_delta_time:units = "seconds since 2018-01-01" ;
  	int end_geoseg(phony_dim_9) ;
  		end_geoseg:contentType = "auxiliaryInformation" ;
  		end_geoseg:description = "The ending geolocation segment number associated with the data contained within this granule. ICESat granule geographic regions are further refined by geolocation segments. During the geolocation process, a geolocation segment is created approximately every 20m from the start of the orbit to the end.  The geolocation segments help align the ATLAS strong a weak beams and provide a common segment length for the L2 and higher products. The geolocation segment indices differ slightly from orbit-to-orbit because of the irregular shape of the Earth. The geolocation segment indices on ATL01 and ATL02 are only approximate because beams have not been aligned at the time of their creation." ;
  		end_geoseg:long_name = "Ending Geolocation Segment" ;
  		end_geoseg:source = "Derived" ;
  		end_geoseg:units = "1" ;
  	double end_gpssow(phony_dim_9) ;
  		end_gpssow:contentType = "auxiliaryInformation" ;
  		end_gpssow:source = "Derived" ;
  		end_gpssow:description = "GPS seconds-of-week of the last data point in the granule." ;
  		end_gpssow:long_name = "Ending GPS SOW of Granule (Actual)" ;
  		end_gpssow:units = "seconds" ;
  	int end_gpsweek(phony_dim_9) ;
  		end_gpsweek:contentType = "auxiliaryInformation" ;
  		end_gpsweek:description = "GPS week number of the last data point in the granule." ;
  		end_gpsweek:long_name = "Ending GPSWeek of Granule (Actual)" ;
  		end_gpsweek:source = "Derived" ;
  		end_gpsweek:units = "weeks from 1980-01-06" ;
  	int end_orbit(phony_dim_9) ;
  		end_orbit:contentType = "auxiliaryInformation" ;
  		end_orbit:description = "The ending orbit number associated with the data contained within this granule. The orbit number increments each time the spacecraft completes a full orbit of the Earth." ;
  		end_orbit:long_name = "Ending Orbit Number" ;
  		end_orbit:source = "Derived" ;
  		end_orbit:units = "1" ;
  	int end_region(phony_dim_9) ;
  		end_region:contentType = "auxiliaryInformation" ;
  		end_region:description = "The ending product-specific region number associated with the data contained within this granule. ICESat-2 data products are separated by geographic regions. The data contained within a specific region are the same for ATL01 and ATL02. ATL03 regions differ slightly because of different geolocation segment locations caused by the irregular shape of the Earth. The region indices for other products are completely independent." ;
  		end_region:long_name = "Ending Region" ;
  		end_region:source = "Derived" ;
  		end_region:units = "1" ;
  	int end_rgt(phony_dim_9) ;
  		end_rgt:contentType = "auxiliaryInformation" ;
  		end_rgt:description = "The ending reference groundtrack (RGT) number associated with the data contained within this granule. There are 1387 reference groundtrack in the ICESat-2 repeat orbit. The reference groundtrack increments each time the spacecraft completes a full orbit of the Earth and resets to 1 each time the spacecraft completes a full cycle." ;
  		end_rgt:long_name = "Ending Reference Groundtrack" ;
  		end_rgt:source = "Derived" ;
  		end_rgt:units = "1" ;
  		end_rgt:valid_max = 1387 ;
  		end_rgt:valid_min = 1 ;
  	string granule_end_utc(phony_dim_9) ;
  		granule_end_utc:contentType = "auxiliaryInformation" ;
  		granule_end_utc:description = "Requested end time (in UTC CCSDS-A) of this granule." ;
  		granule_end_utc:long_name = "End UTC Time of Granule (CCSDS-A, Requested)" ;
  		granule_end_utc:source = "Derived" ;
  		granule_end_utc:units = "1" ;
  	string granule_start_utc(phony_dim_9) ;
  		granule_start_utc:contentType = "auxiliaryInformation" ;
  		granule_start_utc:description = "Requested start time (in UTC CCSDS-A) of this granule." ;
  		granule_start_utc:long_name = "Start UTC Time of Granule (CCSDS-A, Requested)" ;
  		granule_start_utc:source = "Derived" ;
  		granule_start_utc:units = "1" ;
  	double qa_at_interval(phony_dim_9) ;
  		qa_at_interval:contentType = "auxiliaryInformation" ;
  		qa_at_interval:description = "Statistics time interval for along-track QA data." ;
  		qa_at_interval:long_name = "QA Along-Track Interval" ;
  		qa_at_interval:source = "control" ;
  		qa_at_interval:units = "1" ;
  	string release(phony_dim_9) ;
  		release:contentType = "auxiliaryInformation" ;
  		release:description = "Release number of the granule. The release number is incremented when the software or ancillary data used to create the granule has been changed." ;
  		release:long_name = "Release Number" ;
  		release:source = "Operations" ;
  		release:units = "1" ;
  	int start_cycle(phony_dim_9) ;
  		start_cycle:contentType = "auxiliaryInformation" ;
  		start_cycle:description = "The starting cycle number associated with the data contained within this granule. The cycle number is the counter of the number of 91-day repeat cycles completed by the mission." ;
  		start_cycle:long_name = "Starting Cycle" ;
  		start_cycle:source = "Derived" ;
  		start_cycle:units = "1" ;
  		start_cycle:valid_max = 99 ;
  		start_cycle:valid_min = 0 ;
  	double start_delta_time(phony_dim_9) ;
  		start_delta_time:contentType = "auxiliaryInformation" ;
  		start_delta_time:description = "Number of GPS seconds since the ATLAS SDP epoch at the first data point in the file. The ATLAS Standard Data Products (SDP) epoch offset is defined within /ancillary_data/atlas_sdp_gps_epoch as the number of GPS seconds between the GPS epoch (1980-01-06T00:00:00.000000Z UTC) and the ATLAS SDP epoch. By adding the offset contained within atlas_sdp_gps_epoch to delta time parameters, the time in gps_seconds relative to the GPS epoch can be computed." ;
  		start_delta_time:long_name = "ATLAS Start Time (Actual)" ;
  		start_delta_time:source = "Derived" ;
  		start_delta_time:standard_name = "time" ;
  		start_delta_time:units = "seconds since 2018-01-01" ;
  	int start_geoseg(phony_dim_9) ;
  		start_geoseg:contentType = "auxiliaryInformation" ;
  		start_geoseg:description = "The starting geolocation segment number associated with the data contained within this granule. ICESat granule geographic regions are further refined by geolocation segments. During the geolocation process, a geolocation segment is created approximately every 20m from the start of the orbit to the end.  The geolocation segments help align the ATLAS strong a weak beams and provide a common segment length for the L2 and higher products. The geolocation segment indices differ slightly from orbit-to-orbit because of the irregular shape of the Earth. The geolocation segment indices on ATL01 and ATL02 are only approximate because beams have not been aligned at the time of their creation." ;
  		start_geoseg:long_name = "Starting Geolocation Segment" ;
  		start_geoseg:source = "Derived" ;
  		start_geoseg:units = "1" ;
  	double start_gpssow(phony_dim_9) ;
  		start_gpssow:contentType = "auxiliaryInformation" ;
  		start_gpssow:description = "GPS seconds-of-week of the first data point in the granule." ;
  		start_gpssow:long_name = "Start GPS SOW of Granule (Actual)" ;
  		start_gpssow:source = "Derived" ;
  		start_gpssow:units = "seconds" ;
  	int start_gpsweek(phony_dim_9) ;
  		start_gpsweek:contentType = "auxiliaryInformation" ;
  		start_gpsweek:description = "GPS week number of the first data point in the granule." ;
  		start_gpsweek:long_name = "Start GPSWeek of Granule (Actual)" ;
  		start_gpsweek:source = "Derived" ;
  		start_gpsweek:units = "weeks from 1980-01-06" ;
  	int start_orbit(phony_dim_9) ;
  		start_orbit:contentType = "auxiliaryInformation" ;
  		start_orbit:description = "The starting orbit number associated with the data contained within this granule. The orbit number increments each time the spacecraft completes a full orbit of the Earth." ;
  		start_orbit:long_name = "Starting Orbit Number" ;
  		start_orbit:source = "Derived" ;
  		start_orbit:units = "1" ;
  	int start_region(phony_dim_9) ;
  		start_region:contentType = "auxiliaryInformation" ;
  		start_region:description = "The starting product-specific region number associated with the data contained within this granule. ICESat-2 data products are separated by geographic regions. The data contained within a specific region are the same for ATL01 and ATL02. ATL03 regions differ slightly because of different geolocation segment locations caused by the irregular shape of the Earth. The region indices for other products are completely independent." ;
  		start_region:long_name = "Starting Region" ;
  		start_region:source = "Derived" ;
  		start_region:units = "1" ;
  	int start_rgt(phony_dim_9) ;
  		start_rgt:contentType = "auxiliaryInformation" ;
  		start_rgt:description = "The starting reference groundtrack (RGT) number associated with the data contained within this granule. There are 1387 reference groundtrack in the ICESat-2 repeat orbit. The reference groundtrack increments each time the spacecraft completes a full orbit of the Earth and resets to 1 each time the spacecraft completes a full cycle." ;
  		start_rgt:long_name = "Starting Reference Groundtrack" ;
  		start_rgt:source = "Derived" ;
  		start_rgt:units = "1" ;
  		start_rgt:valid_max = 1387 ;
  		start_rgt:valid_min = 1 ;
  	string version(phony_dim_9) ;
  		version:contentType = "auxiliaryInformation" ;
  		version:description = "Version number of this granule within the release. It is a sequential number corresponding to the number of times the granule has been reprocessed for the current release." ;
  		version:long_name = "Version" ;
  		version:source = "Operations" ;
  		version:units = "1" ;

  // group attributes:
  		:Description = "Contains information ancillary to the data product. This may include product characteristics, instrument characteristics and/or processing constants." ;
  		:data_rate = "Data within this group pertain to the granule in its entirety." ;

  group: land {
    dimensions:
    	phony_dim_7 = UNLIMITED ; // (1 currently)
    	phony_dim_8 = 1 ;
    variables:
    	int atl08_region(phony_dim_7) ;
    		atl08_region:contentType = "modelResult" ;
    		atl08_region:description = "ATL08 region(s) encompassed by ATL03 granule being processed" ;
    		atl08_region:long_name = "atl08 region" ;
    		atl08_region:source = "Land ATBD 29March2019, Table 2.4" ;
    		atl08_region:standard_name = "atl08_region" ;
    		atl08_region:units = "1" ;
    	float bin_size_h(phony_dim_8) ;
    		bin_size_h:contentType = "auxiliaryInformation" ;
    		bin_size_h:description = "Histogram bin size for the alternative DRAGANN algorithm. (Default = 1.0)" ;
    		bin_size_h:long_name = "neighbor histogram bin size" ;
    		bin_size_h:source = "ATBD (section 4.2.1 step 3)" ;
    		bin_size_h:units = "1" ;
    	int bin_size_n(phony_dim_8) ;
    		bin_size_n:contentType = "auxiliaryInformation" ;
    		bin_size_n:description = "Size of neighbor histogram bins in number of neighbors in DRAGANN. (Default = 1)" ;
    		bin_size_n:long_name = "neighbor histogram bin size" ;
    		bin_size_n:source = "ATBD (section 4.2 step 4)" ;
    		bin_size_n:units = "1" ;
    	float bright_thresh(phony_dim_8) ;
    		bright_thresh:contentType = "auxiliaryInformation" ;
    		bright_thresh:description = "Threshold to set brightness_flag, average ground photons per shot. (Default = 3.0)" ;
    		bright_thresh:long_name = "brightness flag average ph per shot" ;
    		bright_thresh:source = "ATBD section 2.4.21" ;
    		bright_thresh:units = "1" ;
    	int ca_class(phony_dim_8) ;
    		ca_class:contentType = "auxiliaryInformation" ;
    		ca_class:units = "1" ;
    		ca_class:description = "Canopy classification flag value. (Default = 2)" ;
    		ca_class:long_name = "Canopy class value" ;
    		ca_class:source = "ATBD section 4.12 step 1" ;
    	int can_noise_thresh(phony_dim_8) ;
    		can_noise_thresh:contentType = "auxiliaryInformation" ;
    		can_noise_thresh:units = "1" ;
    		can_noise_thresh:description = "Threshold, as a number of canopy photons in the CAN_FILT_SEG, used for the reclassification of canopy signal photons. (Default = 75)" ;
    		can_noise_thresh:long_name = "Threshold for reclassification of canopy as noise" ;
    		can_noise_thresh:source = "ATBD section 4.11 step 6" ;
    	float can_stat_thresh(phony_dim_8) ;
    		can_stat_thresh:contentType = "auxiliaryInformation" ;
    		can_stat_thresh:units = "1" ;
    		can_stat_thresh:description = "Minimum percentage of canopy photons to compute statistics upon. (Default =0.05)" ;
    		can_stat_thresh:long_name = "Threshold for canopy statistics" ;
    		can_stat_thresh:source = "ATBD section 4.14.1 step 1" ;
    	int canopy_flag_switch(phony_dim_8) ;
    		canopy_flag_switch:contentType = "auxiliaryInformation" ;
    		canopy_flag_switch:source = "ATBD section 4.3" ;
    		canopy_flag_switch:description = "Controls entrance to the canopy flag subroutine . (Default = 1)" ;
    		canopy_flag_switch:long_name = "canopy_flag switch" ;
    		canopy_flag_switch:units = "1" ;
    	int canopy_seg(phony_dim_8) ;
    		canopy_seg:contentType = "auxiliaryInformation" ;
    		canopy_seg:units = "1" ;
    		canopy_seg:description = "Segment in number of signal photons for filtering sparse canopy cover. (Default = 500)" ;
    		canopy_seg:long_name = "segment size in canopy filter" ;
    		canopy_seg:source = "ATBD section 4.11 step 6" ;
    	int class_thresh(phony_dim_8) ;
    		class_thresh:contentType = "auxiliaryInformation" ;
    		class_thresh:description = "Threshold flag value for classification of photons as signal via input from ATL03. (Default =3)" ;
    		class_thresh:long_name = "Threshold flag value for classification of photons as signal via input from ATL03" ;
    		class_thresh:source = "ATBD section 4.2 step 17" ;
    		class_thresh:units = "1" ;
    	int cloud_filter_switch(phony_dim_8) ;
    		cloud_filter_switch:contentType = "auxiliaryInformation" ;
    		cloud_filter_switch:description = "Controls entrance to the cloud_filter subroutine. (Default = 0)" ;
    		cloud_filter_switch:long_name = "cloud_filter switch" ;
    		cloud_filter_switch:source = "ATBD section 4.1.1" ;
    		cloud_filter_switch:units = "1" ;
    	float del_amp(phony_dim_8) ;
    		del_amp:contentType = "auxiliaryInformation" ;
    		del_amp:description = "Step size for optimizing the amplitude variable of Gaussian function. (Default = 1.0)" ;
    		del_amp:long_name = "Step Gaussian Amplitude optimization" ;
    		del_amp:source = "ATBD section 4.2 step 7" ;
    		del_amp:units = "1" ;
    	float del_mu(phony_dim_8) ;
    		del_mu:contentType = "auxiliaryInformation" ;
    		del_mu:description = "Step size for optimizing the mean parameter of Gaussian function. (Default = 0.2)" ;
    		del_mu:long_name = "Step size for optimizing the mean parameter of Gaussian function." ;
    		del_mu:source = "ATBD section 4.2 step 7" ;
    		del_mu:units = "1" ;
    	float del_sigma(phony_dim_8) ;
    		del_sigma:contentType = "auxiliaryInformation" ;
    		del_sigma:description = "Step size for optimizing the standard deviation parameter of Gaussian function. (Default = 0.5)" ;
    		del_sigma:long_name = "Step size for optimizing the standard deviation parameter of Gaussian function." ;
    		del_sigma:source = "ATBD section 4.2 step 7" ;
    		del_sigma:units = "1" ;
    	int dem_filter_switch(phony_dim_8) ;
    		dem_filter_switch:contentType = "auxiliaryInformation" ;
    		dem_filter_switch:description = "Controls filtering based on DEM. (Default = 1)" ;
    		dem_filter_switch:long_name = "dem_filter switch" ;
    		dem_filter_switch:source = "ATBD section 4.5 step 5" ;
    		dem_filter_switch:units = "1" ;
    	float dem_removal_percent_limit(phony_dim_8) ;
    		dem_removal_percent_limit:contentType = "auxiliaryInformation" ;
    		dem_removal_percent_limit:description = "Percent of photons in land segment failing DEM test to set dem_removal_flag. (default = 20.0)" ;
    		dem_removal_percent_limit:long_name = "dem_removal_flag set threshold" ;
    		dem_removal_percent_limit:source = "ATBD section 2.4.11" ;
    		dem_removal_percent_limit:units = "percent" ;
    	int dragann_switch(phony_dim_8) ;
    		dragann_switch:contentType = "auxiliaryInformation" ;
    		dragann_switch:description = "Controls entrance to the DRAGANN subroutine. (Default =1)" ;
    		dragann_switch:long_name = "DRAGANN switch" ;
    		dragann_switch:source = "ATBD section 4.2" ;
    		dragann_switch:units = "1" ;
    	int dseg(phony_dim_8) ;
    		dseg:contentType = "auxiliaryInformation" ;
    		dseg:description = "DRAGANN segment length in 20m geolocated segments along ground track. (Default=170)" ;
    		dseg:long_name = "DRAGANN segment size" ;
    		dseg:source = "ATBD section 4.2.1 step 1" ;
    		dseg:units = "1" ;
    	int dseg_buf(phony_dim_8) ;
    		dseg_buf:contentType = "auxiliaryInformation" ;
    		dseg_buf:description = "DRAGANN segment buffer length in 20m geolocated segments along ground track. (Default=10)" ;
    		dseg_buf:long_name = "DRAGANN segment buffer size" ;
    		dseg_buf:source = "ATBD section 4.2.1 step 1" ;
    		dseg_buf:units = "1" ;
    	int fnlgnd_filter_switch(phony_dim_8) ;
    		fnlgnd_filter_switch:contentType = "auxiliaryInformation" ;
    		fnlgnd_filter_switch:description = "Controls filtering based on FINALGROUND. (Default = 1)" ;
    		fnlgnd_filter_switch:long_name = "finalground filter switch" ;
    		fnlgnd_filter_switch:source = "ATBD section 4.13 step 2" ;
    		fnlgnd_filter_switch:units = "1" ;
    	float gnd_stat_thresh(phony_dim_8) ;
    		gnd_stat_thresh:contentType = "auxiliaryInformation" ;
    		gnd_stat_thresh:description = "Minimum percentage of terrain photons to compute statistics upon. (Default =0.05)" ;
    		gnd_stat_thresh:long_name = "Threshold for terrain statistics" ;
    		gnd_stat_thresh:source = "ATBD section 4.13 step 2" ;
    		gnd_stat_thresh:units = "1" ;
    	float gthresh_factor(phony_dim_8) ;
    		gthresh_factor:contentType = "auxiliaryInformation" ;
    		gthresh_factor:description = "Controls threshold for Gaussian Elimination. (Default = 0.1)" ;
    		gthresh_factor:long_name = "threshold for Gaussian Elimination" ;
    		gthresh_factor:source = "ATBD sGaussian Rejection section of Appendix A" ;
    		gthresh_factor:units = "1" ;
    	float h_canopy_perc(phony_dim_8) ;
    		h_canopy_perc:contentType = "auxiliaryInformation" ;
    		h_canopy_perc:description = "Percentile component of h_canopy parameter. (Default =0.95)" ;
    		h_canopy_perc:long_name = "h_canopy percentile" ;
    		h_canopy_perc:source = "ATBD section 2.2.3" ;
    		h_canopy_perc:units = "1" ;
    	int iter_gnd(phony_dim_8) ;
    		iter_gnd:contentType = "auxiliaryInformation" ;
    		iter_gnd:description = "Iterations of smoothing of interpolated ground surface for refinement. (Default = 10)" ;
    		iter_gnd:long_name = "Iterations of smoothing of interpolated ground surface for ground estimate." ;
    		iter_gnd:source = "ATBD section 4.10 step 1" ;
    		iter_gnd:units = "1" ;
    	int iter_max(phony_dim_8) ;
    		iter_max:contentType = "auxiliaryInformation" ;
    		iter_max:description = "Maximum number of iterations for optimizing the Gaussian parameters for fitting of histogram. (Default = 10)" ;
    		iter_max:long_name = "Maximum number of iterations for optimizing the Gaussian parameters for fitting of histogram." ;
    		iter_max:source = "ATBD section 4.2 step 7" ;
    		iter_max:units = "1" ;
    	int lseg(phony_dim_8) ;
    		lseg:contentType = "auxiliaryInformation" ;
    		lseg:description = "Long segment size in number of 20 meter segments along ground track. (Default=500)" ;
    		lseg:long_name = "Long segment size" ;
    		lseg:source = "ATBD section 4.1 step 1" ;
    		lseg:units = "1" ;
    	int lseg_buf(phony_dim_8) ;
    		lseg_buf:contentType = "auxiliaryInformation" ;
    		lseg_buf:description = "Overlapping long segment buffer size in 20m geosegments along ground track. (Default=10)" ;
    		lseg_buf:long_name = "Long segment buffer size" ;
    		lseg_buf:source = "ATBD section 4.1 step 2" ;
    		lseg_buf:units = "1" ;
    	int lw_filt_bnd(phony_dim_8) ;
    		lw_filt_bnd:contentType = "auxiliaryInformation" ;
    		lw_filt_bnd:description = "Lower bound of the filter window size function. (Default = 5)" ;
    		lw_filt_bnd:long_name = "Proportionality coefficient for controlling the bounds of the filter window size as a function of number of signal photons." ;
    		lw_filt_bnd:source = "ATBD section 4.4 step 2" ;
    		lw_filt_bnd:units = "1" ;
    	float lw_gnd_bnd(phony_dim_8) ;
    		lw_gnd_bnd:contentType = "auxiliaryInformation" ;
    		lw_gnd_bnd:description = "Lower bound restricting the search of a ground surface in canopy cases. (Default = -4.0)" ;
    		lw_gnd_bnd:long_name = "Lower bound restricting the search of a ground surface in canopy cases." ;
    		lw_gnd_bnd:source = "ATBD section 4.7 step 3" ;
    		lw_gnd_bnd:units = "meters" ;
    	float lw_toc_bnd(phony_dim_8) ;
    		lw_toc_bnd:contentType = "auxiliaryInformation" ;
    		lw_toc_bnd:description = "Lower bound restricting the search of a top of canopy surface. (Default = -4.0)" ;
    		lw_toc_bnd:long_name = "Lower bound restricting the search of a top of canopy surface." ;
    		lw_toc_bnd:source = "section 4.7 step 3 entered from section 4.8" ;
    		lw_toc_bnd:units = "meters" ;
    	float lw_toc_cut(phony_dim_8) ;
    		lw_toc_cut:contentType = "auxiliaryInformation" ;
    		lw_toc_cut:description = "Lower cutoff for top of canopy surface. (Default = 2.0)" ;
    		lw_toc_cut:long_name = "Lower cutoff for top of canopy" ;
    		lw_toc_cut:source = "ATBD section 4.8 step 10" ;
    		lw_toc_cut:units = "meters" ;
    	int max_atl03files(phony_dim_8) ;
    		max_atl03files:contentType = "auxiliaryInformation" ;
    		max_atl03files:description = "Maximum number of input ATL03 files. (Default = 200)" ;
    		max_atl03files:long_name = "Maximum number of input ATL03s" ;
    		max_atl03files:source = "Operations" ;
    		max_atl03files:units = "1" ;
    	int max_atl09files(phony_dim_8) ;
    		max_atl09files:contentType = "auxiliaryInformation" ;
    		max_atl09files:description = "Maximum number of input ATL09 files. (Default = 200)" ;
    		max_atl09files:long_name = "Maximum number of input ATL09s" ;
    		max_atl09files:source = "Operations" ;
    		max_atl09files:units = "1" ;
    	int max_peaks(phony_dim_8) ;
    		max_peaks:contentType = "auxiliaryInformation" ;
    		max_peaks:source = "ATBD section 4.2 step 9" ;
    		max_peaks:description = "Maximum number of Gaussian peaks to fit in the data set in DRAGANN. (Default =10)" ;
    		max_peaks:long_name = "Maximum number of Gaussian peaks to fit in the data set" ;
    		max_peaks:units = "1" ;
    	int max_try(phony_dim_8) ;
    		max_try:contentType = "auxiliaryInformation" ;
    		max_try:description = "Maximum number of tries to compute a P value in alternative DRAGANN" ;
    		max_try:long_name = "Maximum try count" ;
    		max_try:source = "ATBD section 4.2.1 step 17" ;
    		max_try:units = "1" ;
    	int min_nphs(phony_dim_8) ;
    		min_nphs:contentType = "auxiliaryInformation" ;
    		min_nphs:description = "Minimum number of input photons from ATL03 to process. (default=1)" ;
    		min_nphs:long_name = "Minimum input photons" ;
    		min_nphs:source = "Operations" ;
    		min_nphs:units = "1" ;
    	int n_dec_mode(phony_dim_8) ;
    		n_dec_mode:contentType = "auxiliaryInformation" ;
    		n_dec_mode:description = "Number of decimal places to consider in mode computation. (Default =1)" ;
    		n_dec_mode:long_name = "Mode decimal parameter" ;
    		n_dec_mode:source = "ATBD needed for section 4.13 step 3(h_te_mode)" ;
    		n_dec_mode:units = "1" ;
    	float night_thresh(phony_dim_8) ;
    		night_thresh:contentType = "auxiliaryInformation" ;
    		night_thresh:description = "Solar elevation threshold for determining night time conditions. (Default =0.0)" ;
    		night_thresh:long_name = "Threshold for night" ;
    		night_thresh:source = "ATBD section 2.4.9" ;
    		night_thresh:units = "1" ;
    	int noise_class(phony_dim_8) ;
    		noise_class:contentType = "auxiliaryInformation" ;
    		noise_class:description = "Noise classification flag value. (Default = 0)" ;
    		noise_class:long_name = "Noise class value" ;
    		noise_class:source = "ATBD section 4.12 step 1" ;
    		noise_class:units = "1" ;
    	int outlier_filter_switch(phony_dim_8) ;
    		outlier_filter_switch:contentType = "auxiliaryInformation" ;
    		outlier_filter_switch:description = "Controls entrance to the outlier filter subroutine. (Default = 1)" ;
    		outlier_filter_switch:long_name = "outlier_filter switch" ;
    		outlier_filter_switch:source = "ATBD section 4.6" ;
    		outlier_filter_switch:units = "1" ;
    	float p_static(phony_dim_8) ;
    		p_static:contentType = "auxiliaryInformation" ;
    		p_static:description = "Parameter for controlling the search radius in nearest neighbor search in DRAGANN. (Default = 20)" ;
    		p_static:long_name = "Dragann Parameter" ;
    		p_static:source = "ATBD section 4.2 step 1" ;
    		p_static:units = "1" ;
    	float ph_removal_percent_limit(phony_dim_8) ;
    		ph_removal_percent_limit:contentType = "auxiliaryInformation" ;
    		ph_removal_percent_limit:description = "Percent of photons in land segment removed to set ph_removal_flag. (default = 50.0)" ;
    		ph_removal_percent_limit:long_name = "ph_removal_flag set threshold" ;
    		ph_removal_percent_limit:source = "ATBD section 4.13 step 4" ;
    		ph_removal_percent_limit:units = "percent" ;
    	int proc_geoseg(phony_dim_8) ;
    		proc_geoseg:contentType = "auxiliaryInformation" ;
    		proc_geoseg:description = "Geosegment process interval length.  This controls the amount read from ATL03 and ATL09 at a time. (Default = 500000)." ;
    		proc_geoseg:long_name = "Geosegment process interval length" ;
    		proc_geoseg:source = "Operations" ;
    		proc_geoseg:units = "1" ;
    	float psf(phony_dim_8) ;
    		psf:contentType = "auxiliaryInformation" ;
    		psf:description = "Parameter controlling identification of photons around an interpolated surface. (Default = 0.5)" ;
    		psf:long_name = "Point Spread Function" ;
    		psf:source = "ATBD section 4.7 step 12" ;
    		psf:units = "meters" ;
    	float ref_dem_limit(phony_dim_8) ;
    		ref_dem_limit:contentType = "auxiliaryInformation" ;
    		ref_dem_limit:description = "Reference DEM limit used to reclassify signal as noise. (default = 120.0)" ;
    		ref_dem_limit:long_name = "DEM threshold" ;
    		ref_dem_limit:source = "ATBD section 4.5 step 4" ;
    		ref_dem_limit:units = "meters" ;
    	float ref_finalground_limit(phony_dim_8) ;
    		ref_finalground_limit:contentType = "auxiliaryInformation" ;
    		ref_finalground_limit:units = "meters" ;
    		ref_finalground_limit:description = "Reference finalground limit used to reclassify signal as noise. (default = 150.0)" ;
    		ref_finalground_limit:long_name = "finalground threshold" ;
    		ref_finalground_limit:source = "ATBD section 4.13 step 2" ;
    	float relief_hbot(phony_dim_8) ;
    		relief_hbot:contentType = "auxiliaryInformation" ;
    		relief_hbot:description = "The approximate relief of the L-km segment uses the percentile height values, relief_htop and relief_hbot. (Default=0.05)" ;
    		relief_hbot:long_name = "lower relief percentile" ;
    		relief_hbot:source = "ATBD (section 4.5 step 6)" ;
    		relief_hbot:units = "meters" ;
    	float relief_htop(phony_dim_8) ;
    		relief_htop:contentType = "auxiliaryInformation" ;
    		relief_htop:description = "The approximate relief of the L-km segment uses the percentile height values, relief_htop and relief_hbot. (Default=0.95)" ;
    		relief_htop:long_name = "Upper relief percentile" ;
    		relief_htop:source = "ATBD (section 4.5 step 6)" ;
    		relief_htop:units = "meters" ;
    	float shp_param(phony_dim_8) ;
    		shp_param:contentType = "auxiliaryInformation" ;
    		shp_param:description = "Exponential coefficient of the filter window size as a function. (Default = 21.0E-06)" ;
    		shp_param:long_name = "Exponential coefficient for controlling the exponential decay of the filter window size as a function of number of signal photons." ;
    		shp_param:source = "ATBD section 4.4 step 2" ;
    		shp_param:units = "1" ;
    	float sig_rsq_search(phony_dim_8) ;
    		sig_rsq_search:contentType = "auxiliaryInformation" ;
    		sig_rsq_search:description = "Top of canopy refinement square search radius. (Default = 225.0)" ;
    		sig_rsq_search:long_name = "Square Radius of filter for canopy" ;
    		sig_rsq_search:source = "ATBD section 4.8 step 6" ;
    		sig_rsq_search:units = "meters^2" ;
    	float sseg(phony_dim_8) ;
    		sseg:contentType = "auxiliaryInformation" ;
    		sseg:description = "Short segment length in meters. (Default = 100.0)" ;
    		sseg:long_name = "Short Segment Length" ;
    		sseg:source = "ATBD section 4.13 step 1" ;
    		sseg:units = "meters" ;
    	int stat_thresh(phony_dim_8) ;
    		stat_thresh:contentType = "auxiliaryInformation" ;
    		stat_thresh:description = "Minimum number of photons to compute statistics upon. (Default =50)" ;
    		stat_thresh:long_name = "Threshold for land statistics" ;
    		stat_thresh:source = "ATBD section 2 intro paragraph" ;
    		stat_thresh:units = "1" ;
    	float tc_thresh(phony_dim_8) ;
    		tc_thresh:contentType = "auxiliaryInformation" ;
    		tc_thresh:description = "Percentage threshold for average L-km segment tree cover to be considered canopy. (Default = 5.0)" ;
    		tc_thresh:long_name = "Canopy Flag threshold" ;
    		tc_thresh:source = "ATBD section 4.3 steps 6 and 7" ;
    		tc_thresh:units = "1" ;
    	int te_class(phony_dim_8) ;
    		te_class:contentType = "auxiliaryInformation" ;
    		te_class:description = "Terrain classification flag value. (Default = 1)" ;
    		te_class:long_name = "Terrain class value" ;
    		te_class:source = "ATBD section 4.12 step 1" ;
    		te_class:units = "1" ;
    	int toc_class(phony_dim_8) ;
    		toc_class:contentType = "auxiliaryInformation" ;
    		toc_class:description = "Top of canopy classification flag value. (Default = 3)" ;
    		toc_class:long_name = "Top of canopy class value" ;
    		toc_class:source = "ATBD section 4.12 step 1" ;
    		toc_class:units = "1" ;
    	int up_filt_bnd(phony_dim_8) ;
    		up_filt_bnd:contentType = "auxiliaryInformation" ;
    		up_filt_bnd:description = "Lower bound of the filter window size function. (Default = 46)" ;
    		up_filt_bnd:long_name = "Proportionality coefficient for controlling the bounds of the filter window size as a function of number of signal photons." ;
    		up_filt_bnd:source = "ATBD section 4.4 step 2" ;
    		up_filt_bnd:units = "1" ;
    	float up_gnd_bnd(phony_dim_8) ;
    		up_gnd_bnd:contentType = "auxiliaryInformation" ;
    		up_gnd_bnd:description = "Upper bound restricting the search of a ground surface in canopy cases. (Default = 1.0)" ;
    		up_gnd_bnd:long_name = "Upper bound restricting the search of a ground surface in canopy cases." ;
    		up_gnd_bnd:source = "ATBD (section 4.7 step 3)" ;
    		up_gnd_bnd:units = "meters" ;
    	float up_toc_bnd(phony_dim_8) ;
    		up_toc_bnd:contentType = "auxiliaryInformation" ;
    		up_toc_bnd:description = "Upper bound restricting the search of a top of canopy surface. (Default=1.0)" ;
    		up_toc_bnd:long_name = "Upper bound restricting the search of a top of canopy surface." ;
    		up_toc_bnd:source = "ATBD section 4.7 step 3 entered from section 4.8" ;
    		up_toc_bnd:units = "meters" ;
    	float up_toc_cut(phony_dim_8) ;
    		up_toc_cut:contentType = "auxiliaryInformation" ;
    		up_toc_cut:description = "Upper cutoff for top of canopy surface. (Default = 150.0)" ;
    		up_toc_cut:long_name = "upper cutoff of top of canopy surface." ;
    		up_toc_cut:source = "ATBD section 4.8 step 10" ;
    		up_toc_cut:units = "meters" ;

    // group attributes:
    		:Description = "Constants used in the land_vegetation ATBD" ;
    } // group land
  } // group ancillary_data

group: orbit_info {
  dimensions:
  	crossing_time = UNLIMITED ; // (1 currently)
  	sc_orient_time = UNLIMITED ; // (1 currently)
  variables:
  	double crossing_time(crossing_time) ;
  		crossing_time:contentType = "referenceInformation" ;
  		crossing_time:description = "The time, in seconds since the ATLAS SDP GPS Epoch, at which the ascending node crosses the equator. The ATLAS Standard Data Products (SDP) epoch offset is defined within /ancillary_data/atlas_sdp_gps_epoch as the number of GPS seconds between the GPS epoch (1980-01-06T00:00:00.000000Z UTC) and the ATLAS SDP epoch. By adding the offset contained within atlas_sdp_gps_epoch to delta time parameters, the time in gps_seconds relative to the GPS epoch can be computed." ;
  		crossing_time:long_name = "Ascending Node Crossing Time" ;
  		crossing_time:source = "POD/PPD" ;
  		crossing_time:standard_name = "time" ;
  		crossing_time:units = "seconds since 2018-01-01" ;
  	byte cycle_number(crossing_time) ;
  		cycle_number:contentType = "referenceInformation" ;
  		cycle_number:coordinates = "crossing_time" ;
  		cycle_number:description = "A count of the number of exact repeats of this reference orbit." ;
  		cycle_number:long_name = "Cycle Number" ;
  		cycle_number:source = "Operations" ;
  		cycle_number:units = "1" ;
  		cycle_number:valid_max = 50b ;
  		cycle_number:valid_min = 0b ;
  	double lan(crossing_time) ;
  		lan:contentType = "referenceInformation" ;
  		lan:coordinates = "crossing_time" ;
  		lan:description = "Longitude at the ascending node crossing." ;
  		lan:long_name = "Ascending Node Longitude" ;
  		lan:source = "POD/PPD" ;
  		lan:units = "degrees_east" ;
  		lan:valid_max = 180. ;
  		lan:valid_min = -180. ;
  	ushort orbit_number(crossing_time) ;
  		orbit_number:contentType = "referenceInformation" ;
  		orbit_number:coordinates = "crossing_time" ;
  		orbit_number:description = "Unique identifying number for each planned ICESat-2 orbit." ;
  		orbit_number:long_name = "Orbit Number" ;
  		orbit_number:source = "Operations" ;
  		orbit_number:units = "1" ;
  		orbit_number:valid_max = 65000US ;
  		orbit_number:valid_min = 1US ;
  	short rgt(crossing_time) ;
  		rgt:contentType = "referenceInformation" ;
  		rgt:coordinates = "crossing_time" ;
  		rgt:description = "The reference ground track (RGT) is the track on the earth at which a specified unit vector within the observatory is pointed. Under nominal operating conditions, there will be no data collected along the RGT, as the RGT is spanned by GT3 and GT4.  During slews or off-pointing, it is possible that ground tracks may intersect the RGT. The ICESat-2 mission has 1387 RGTs." ;
  		rgt:long_name = "Reference Ground track" ;
  		rgt:source = "POD/PPD" ;
  		rgt:units = "1" ;
  		rgt:valid_max = 1387s ;
  		rgt:valid_min = 1s ;
  	byte sc_orient(sc_orient_time) ;
  		sc_orient:contentType = "referenceInformation" ;
  		sc_orient:coordinates = "sc_orient_time" ;
  		sc_orient:description = "This parameter tracks the spacecraft orientation between forward, backward and transitional flight modes. ICESat-2 is considered to be flying forward when the weak beams are leading the strong beams; and backward when the strong beams are leading the weak beams. ICESat-2 is considered to be in transition while it is maneuvering between the two orientations. Science quality is potentially degraded while in transition mode." ;
  		sc_orient:flag_meanings = "backward forward transition" ;
  		sc_orient:flag_values = 0b, 1b, 2b ;
  		sc_orient:long_name = "Spacecraft Orientation" ;
  		sc_orient:source = "POD/PPD" ;
  		sc_orient:units = "1" ;
  		sc_orient:valid_max = 2b ;
  		sc_orient:valid_min = 0b ;
  	double sc_orient_time(sc_orient_time) ;
  		sc_orient_time:contentType = "referenceInformation" ;
  		sc_orient_time:description = "The time of the last spacecraft orientation change between forward, backward and transitional flight modes, expressed in seconds since the ATLAS SDP GPS Epoch. ICESat-2 is considered to be flying forward when the weak beams are leading the strong beams; and backward when the strong beams are leading the weak beams. ICESat-2 is considered to be in transition while it is maneuvering between the two orientations. Science quality is potentially degraded while in transition mode. The ATLAS Standard Data Products (SDP) epoch offset is defined within /ancillary_data/atlas_sdp_gps_epoch as the number of GPS seconds between the GPS epoch (1980-01-06T00:00:00.000000Z UTC) and the ATLAS SDP epoch. By adding the offset contained within atlas_sdp_gps_epoch to delta time parameters, the time in gps_seconds relative to the GPS epoch can be computed." ;
  		sc_orient_time:long_name = "Time of Last Spacecraft Orientation Change" ;
  		sc_orient_time:source = "POD/PPD" ;
  		sc_orient_time:standard_name = "time" ;
  		sc_orient_time:units = "seconds since 2018-01-01" ;

  // group attributes:
  		:Description = "Contains orbit information." ;
  		:data_rate = "Varies. Data are only provided when one of the stored values (besides time) changes." ;
  } // group orbit_info

group: quality_assessment {
  dimensions:
  	phony_dim_10 = 1 ;
  variables:
  	int qa_granule_fail_reason(phony_dim_10) ;
  		qa_granule_fail_reason:contentType = "qualityInformation" ;
  		qa_granule_fail_reason:description = "Flag indicating granule failure reason. 0=no failure; 1=processing error; 2=Insufficient output data was generated; 3=TBD Failure; 4=TBD_Failure; 5=other failure." ;
  		qa_granule_fail_reason:flag_meanings = "no_failure PROCESS_ERROR INSUFFICIENT_OUTPUT failure_3 failure_4 OTHER_FAILURE" ;
  		qa_granule_fail_reason:flag_values = 0, 1, 2, 3, 4, 5 ;
  		qa_granule_fail_reason:long_name = "Granule Failure Reason" ;
  		qa_granule_fail_reason:source = "Operations" ;
  		qa_granule_fail_reason:units = "1" ;
  		qa_granule_fail_reason:valid_max = 5 ;
  		qa_granule_fail_reason:valid_min = 0 ;
  	int qa_granule_pass_fail(phony_dim_10) ;
  		qa_granule_pass_fail:contentType = "qualityInformation" ;
  		qa_granule_pass_fail:description = "Flag indicating granule quality. 0=granule passes automatic QA. 1=granule fails automatic QA." ;
  		qa_granule_pass_fail:flag_meanings = "PASS FAIL" ;
  		qa_granule_pass_fail:flag_values = 0, 1 ;
  		qa_granule_pass_fail:long_name = "Granule Pass Flag" ;
  		qa_granule_pass_fail:source = "Operations" ;
  		qa_granule_pass_fail:units = "1" ;
  		qa_granule_pass_fail:valid_max = 1 ;
  		qa_granule_pass_fail:valid_min = 0 ;

  // group attributes:
  		:Description = "Contains quality assessment data. This may include QA counters, QA along-track data and/or QA summary data." ;
  } // group quality_assessment

group: METADATA {

  // group attributes:
  		:Description = "ISO19115 Structured Metadata Represented within HDF5" ;
  		:iso_19139_dataset_xml = "<?xml version=\"1.0\"?>\n<gmd:DS_Series xsi:schemaLocation=\"http://www.isotc211.org/2005/gmi http://cdn.earthdata.nasa.gov/iso/schema/1.0/ISO19115-2_EOS.xsd\" xmlns:eos=\"http://earthdata.nasa.gov/schema/eos\" xmlns:gco=\"http://www.isotc211.org/2005/gco\" xmlns:gmd=\"http://www.isotc211.org/2005/gmd\" xmlns:gmi=\"http://www.isotc211.org/2005/gmi\" xmlns:gml=\"http://www.opengis.net/gml/3.2\" xmlns:gmx=\"http://www.isotc211.org/2005/gmx\" xmlns:gsr=\"http://www.isotc211.org/2005/gsr\" xmlns:gss=\"http://www.isotc211.org/2005/gss\" xmlns:gts=\"http://www.isotc211.org/2005/gts\" xmlns:srv=\"http://www.isotc211.org/2005/srv\" xmlns:xlink=\"http://www.w3.org/1999/xlink\" xmlns:xs=\"http://www.w3.org/2001/XMLSchema\" xmlns:xsi=\"http://www.w3.org/2001/XMLSchema-instance\">\n  <gmd:composedOf>\n    <gmd:DS_DataSet>\n      <gmd:has>\n        <gmi:MI_Metadata>\n          <gmd:fileIdentifier>\n            <gmx:FileName>ATL08_20181014084920_02400109_003_01.h5</gmx:FileName>\n          </gmd:fileIdentifier>\n          <gmd:contact>\n            <gmd:CI_ResponsibleParty>\n              <gmd:organisationName>\n                <gco:CharacterString>NSIDC DAAC &gt; National Snow and Ice Data Center DAAC</gco:CharacterString>\n              </gmd:organisationName>\n              <gmd:contactInfo>\n                <gmd:CI_Contact>\n                  <gmd:address>\n                    <gmd:CI_Address>\n                      <gmd:electronicMailAddress>\n                        <gco:CharacterString>nsidc@nsidc.org</gco:CharacterString>\n                      </gmd:electronicMailAddress>\n                    </gmd:CI_Address>\n                  </gmd:address>\n                  <gmd:onlineResource>\n                    <gmd:CI_OnlineResource>\n                      <gmd:linkage>\n                        <gmd:URL>http://nsidc.org/daac/</gmd:URL>\n                      </gmd:linkage>\n                    </gmd:CI_OnlineResource>\n                  </gmd:onlineResource>\n                </gmd:CI_Contact>\n              </gmd:contactInfo>\n              <gmd:role>\n                <gmd:CI_RoleCode codeList=\"http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_RoleCode\" codeListValue=\"pointOfContact\">pointOfContact</gmd:CI_RoleCode>\n              </gmd:role>\n            </gmd:CI_ResponsibleParty>\n          </gmd:contact>\n          <gmd:dateStamp>\n            <gco:DateTime>2020-04-01T14:03:26.000000Z</gco:DateTime>\n          </gmd:dateStamp>\n          <gmd:identificationInfo>\n            <gmd:MD_DataIdentification>\n              <gmd:citation>\n                <gmd:CI_Citation>\n                  <gmd:title>\n                    <gmx:FileName>ATL08_20181014084920_02400109_003_01.h5</gmx:FileName>\n                  </gmd:title>\n                  <gmd:date>\n                    <gmd:CI_Date>\n                      <gmd:date>\n                        <gco:DateTime>2020-04-01T14:03:26.000000Z</gco:DateTime>\n                      </gmd:date>\n                      <gmd:dateType>\n                        <gmd:CI_DateTypeCode codeList=\"http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode\" codeListValue=\"creation\">creation</gmd:CI_DateTypeCode>\n                      </gmd:dateType>\n                    </gmd:CI_Date>\n                  </gmd:date>\n                  <gmd:identifier>\n                    <gmd:MD_Identifier>\n                      <gmd:code>\n                        <gco:CharacterString>ATL08</gco:CharacterString>\n                      </gmd:code>\n                      <gmd:description>\n                        <gco:CharacterString>The ECS Short Name</gco:CharacterString>\n                      </gmd:description>\n                    </gmd:MD_Identifier>\n                  </gmd:identifier>\n                  <gmd:identifier>\n                    <gmd:MD_Identifier>\n                      <gmd:code>\n                        <gco:CharacterString>003</gco:CharacterString>\n                      </gmd:code>\n                      <gmd:description>\n                        <gco:CharacterString>The ECS Version ID</gco:CharacterString>\n                      </gmd:description>\n                    </gmd:MD_Identifier>\n                  </gmd:identifier>\n                  <gmd:identifier>\n                    <gmd:MD_Identifier>\n                      <gmd:code>\n                        <gco:CharacterString>ATL08_20181014084920_02400109_003_01.h5</gco:CharacterString>\n                      </gmd:code>\n                      <gmd:description>\n                        <gco:CharacterString>ProducerGranuleId</gco:CharacterString>\n                      </gmd:description>\n                    </gmd:MD_Identifier>\n                  </gmd:identifier>\n                </gmd:CI_Citation>\n              </gmd:citation>\n              <gmd:abstract>\n                <gco:CharacterString>The ICESat-2 ATL08 standard data product contains along-track heights of ground and canopy surface at varying length scales. Where data permits, this includes estimates of canopy height, relative canopy cover, canopy height distributions, surface roughness, surface slope/aspect, and apparent reflectance.</gco:CharacterString>\n              </gmd:abstract>\n              <gmd:aggregationInfo>\n                <gmd:MD_AggregateInformation>\n                  <gmd:aggregateDataSetName>\n                    <gmd:CI_Citation>\n                      <gmd:title>\n                        <gco:CharacterString>ATL08</gco:CharacterString>\n                      </gmd:title>\n                      <gmd:date gco:nilReason=\"unknown\"/>\n                      <gmd:edition>\n                        <gco:CharacterString>003</gco:CharacterString>\n                      </gmd:edition>\n                    </gmd:CI_Citation>\n                  </gmd:aggregateDataSetName>\n                  <gmd:associationType>\n                    <gmd:DS_AssociationTypeCode codeList=\"http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#DS_AssociationTypeCode\" codeListValue=\"largerWorkCitation\">largerWorkCitation</gmd:DS_AssociationTypeCode>\n                  </gmd:associationType>\n                </gmd:MD_AggregateInformation>\n              </gmd:aggregationInfo>\n              <gmd:language>\n                <gco:CharacterString>eng</gco:CharacterString>\n              </gmd:language>\n             <gmd:extent>\n                <gmd:EX_Extent id=\"boundingExtent\">\n                  <gmd:geographicElement>\n                    <gmd:EX_GeographicDescription id=\"Orbit\">\n                      <gmd:geographicIdentifier>\n                        <gmd:MD_Identifier>\n                          <gmd:code>\n                            <gco:CharacterString>AscendingCrossing: 114.85413503237267 StartLatitude: -27.000000000000000 StartDirection:D EndLatitude: -50.000000000000000 EndDirection: D</gco:CharacterString>\n                          </gmd:code>\n                          <gmd:codeSpace>\n                            <gco:CharacterString>gov.nasa.esdis.umm.orbitparameters</gco:CharacterString>\n                          </gmd:codeSpace>\n                          <gmd:description>\n                            <gco:CharacterString>OrbitParameters</gco:CharacterString>\n                          </gmd:description>\n                        </gmd:MD_Identifier>\n                      </gmd:geographicIdentifier>\n                    </gmd:EX_GeographicDescription>\n                  </gmd:geographicElement>\n                  <gmd:geographicElement>\n                    <gmd:EX_GeographicDescription id=\"OrbitCalculatedSpatialDomains0\">\n                      <gmd:geographicIdentifier>\n                        <gmd:MD_Identifier>\n                          <gmd:code>\n                            <gco:CharacterString>OrbitNumber: 441 EquatorCrossingLongitude: 114.85413503237267 EquatorCrossingDateTime: 2018-10-14T07:55:13.897432Z</gco:CharacterString>\n                          </gmd:code>\n                          <gmd:codeSpace>\n                            <gco:CharacterString>gov.nasa.esdis.umm.orbitcalculatedspatialdomains</gco:CharacterString>\n                          </gmd:codeSpace>\n                          <gmd:description>\n                            <gco:CharacterString>OrbitCalculatedSpatialDomains</gco:CharacterString>\n                          </gmd:description>\n                        </gmd:MD_Identifier>\n                      </gmd:geographicIdentifier>\n                    </gmd:EX_GeographicDescription>\n                  </gmd:geographicElement>\n                  <gmd:temporalElement>\n                    <gmd:EX_TemporalExtent>\n                      <gmd:extent>\n                        <gml:TimePeriod gml:id=\"TIME_PERIOD_ID\">\n                          <gml:beginPosition>2018-10-14T08:51:05.104949Z</gml:beginPosition>\n                          <gml:endPosition>2018-10-14T08:51:05.172649Z</gml:endPosition>\n                        </gml:TimePeriod>\n                      </gmd:extent>\n                    </gmd:EX_TemporalExtent>\n                  </gmd:temporalElement>\n                </gmd:EX_Extent>\n              </gmd:extent>\n            </gmd:MD_DataIdentification>\n          </gmd:identificationInfo>\n          <gmd:dataQualityInfo>\n            <gmd:DQ_DataQuality>\n              <gmd:scope>\n                <gmd:DQ_Scope>\n                  <gmd:level>\n                    <gmd:MD_ScopeCode codeList=\"http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_ScopeCode\" codeListValue=\"dataset\">dataset</gmd:MD_ScopeCode>\n                  </gmd:level>\n                </gmd:DQ_Scope>\n              </gmd:scope>\n              <gmd:lineage>\n                <gmd:LI_Lineage>\n                  <gmd:processStep>\n                    <gmi:LE_ProcessStep>\n                      <gmd:description>\n                        <gco:CharacterString>2020-04-01T14:03:26.000000Z;ae899cbd-cf20-3541-9952-cb5220d5467b;Created by PGE atlas_l3a_ld Version 3.3.1</gco:CharacterString>\n                      </gmd:description>\n                      <gmd:dateTime>\n                        <gco:DateTime>2020-04-01T14:03:26.000000Z</gco:DateTime>\n                      </gmd:dateTime>\n                    </gmi:LE_ProcessStep>\n                  </gmd:processStep>\n                </gmd:LI_Lineage>\n              </gmd:lineage>\n            </gmd:DQ_DataQuality>\n          </gmd:dataQualityInfo>\n        </gmi:MI_Metadata>\n      </gmd:has>\n    </gmd:DS_DataSet>\n  </gmd:composedOf>\n  <gmd:seriesMetadata gco:nilReason=\"missing\"/>\n</gmd:DS_Series>\n" ;
  		:iso_19139_series_xml = "<?xml version=\"1.0\" encoding=\"UTF-8\"?>\r\n<gmd:DS_Series\r\n  xmlns:eos=\"http://earthdata.nasa.gov/schema/eos\"\r\n  xmlns:gco=\"http://www.isotc211.org/2005/gco\"\r\n  xmlns:gmd=\"http://www.isotc211.org/2005/gmd\"\r\n  xmlns:gmi=\"http://www.isotc211.org/2005/gmi\"\r\n  xmlns:gml=\"http://www.opengis.net/gml/3.2\"\r\n  xmlns:gmx=\"http://www.isotc211.org/2005/gmx\"\r\n  xmlns:gsr=\"http://www.isotc211.org/2005/gsr\"\r\n  xmlns:gss=\"http://www.isotc211.org/2005/gss\"\r\n  xmlns:gts=\"http://www.isotc211.org/2005/gts\"\r\n  xmlns:srv=\"http://www.isotc211.org/2005/srv\"\r\n  xmlns:xlink=\"http://www.w3.org/1999/xlink\"\r\n  xmlns:xs=\"http://www.w3.org/2001/XMLSchema\"\r\n  xmlns:xsi=\"http://www.w3.org/2001/XMLSchema-instance\"\r\n  xsi:schemaLocation=\"http://www.isotc211.org/2005/gmi http://cdn.earthdata.nasa.gov/iso/schema/1.0/ISO19115-2_EOS.xsd\">\r\n  <gmd:composedOf gco:nilReason=\"inapplicable\"/>\r\n  <gmd:seriesMetadata>\r\n    <gmi:MI_Metadata>\r\n      <gmd:fileIdentifier>\r\n        <gco:CharacterString>ATL08.003</gco:CharacterString>\r\n      </gmd:fileIdentifier>\r\n      <gmd:language>\r\n        <gco:CharacterString>eng</gco:CharacterString>\r\n      </gmd:language>\r\n      <gmd:characterSet>\r\n        <gmd:MD_CharacterSetCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#MD_CharacterSetCode\" codeListValue=\"utf8\">utf8</gmd:MD_CharacterSetCode>\r\n      </gmd:characterSet>\r\n      <gmd:hierarchyLevel>\r\n        <gmd:MD_ScopeCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#MD_ScopeCode\" codeListValue=\"series\">series</gmd:MD_ScopeCode>\r\n      </gmd:hierarchyLevel>\r\n      <gmd:contact>\r\n        <gmd:CI_ResponsibleParty>\r\n          <gmd:organisationName>\r\n            <gco:CharacterString>NSIDC DAAC &gt; NASA National Snow and Ice Data Center Distributed Active Archive Center</gco:CharacterString>\r\n          </gmd:organisationName>\r\n          <gmd:contactInfo>\r\n            <gmd:CI_Contact id=\"NSIDC_DAAC_CONTACT_ID\">\r\n              <gmd:phone>\r\n                <gmd:CI_Telephone>\r\n                  <gmd:voice>\r\n                    <gco:CharacterString>303-492-6199</gco:CharacterString>\r\n                  </gmd:voice>\r\n                  <gmd:facsimile>\r\n                    <gco:CharacterString>303-492-2468</gco:CharacterString>\r\n                  </gmd:facsimile>\r\n                </gmd:CI_Telephone>\r\n              </gmd:phone>\r\n              <gmd:address>\r\n                <gmd:CI_Address>\r\n                  <gmd:deliveryPoint>\r\n                    <gco:CharacterString>1540 30th St Campus Box 449</gco:CharacterString>\r\n                  </gmd:deliveryPoint>\r\n                  <gmd:city>\r\n                    <gco:CharacterString>Boulder</gco:CharacterString>\r\n                  </gmd:city>\r\n                  <gmd:administrativeArea>\r\n                    <gco:CharacterString>Colorado</gco:CharacterString>\r\n                  </gmd:administrativeArea>\r\n                  <gmd:postalCode>\r\n                    <gco:CharacterString>80309-0449</gco:CharacterString>\r\n                  </gmd:postalCode>\r\n                  <gmd:country>\r\n                    <gco:CharacterString>USA</gco:CharacterString>\r\n                  </gmd:country>\r\n                  <gmd:electronicMailAddress>\r\n                    <gco:CharacterString>nsidc@nsidc.org</gco:CharacterString>\r\n                  </gmd:electronicMailAddress>\r\n                </gmd:CI_Address>\r\n              </gmd:address>\r\n              <gmd:onlineResource>\r\n                <gmd:CI_OnlineResource>\r\n                  <gmd:linkage>\r\n                    <gmd:URL>http://nsidc.org/daac/</gmd:URL>\r\n                  </gmd:linkage>\r\n                </gmd:CI_OnlineResource>\r\n              </gmd:onlineResource>\r\n              <gmd:hoursOfService>\r\n                <gco:CharacterString>9:00 A.M. to 5:00 P.M., U.S. Mountain Time, Monday through Friday, excluding U.S. holidays.</gco:CharacterString>\r\n              </gmd:hoursOfService>\r\n              <gmd:contactInstructions>\r\n                <gco:CharacterString>Contact by e-mail first</gco:CharacterString>\r\n              </gmd:contactInstructions>\r\n            </gmd:CI_Contact>\r\n          </gmd:contactInfo>\r\n          <gmd:role>\r\n            <gmd:CI_RoleCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#CI_RoleCode\" codeListValue=\"pointOfContact\">pointOfContact</gmd:CI_RoleCode>\r\n          </gmd:role>\r\n        </gmd:CI_ResponsibleParty>\r\n      </gmd:contact>\r\n      <gmd:dateStamp>\r\n        <gco:Date>2015-10-15</gco:Date>\r\n      </gmd:dateStamp>\r\n      <gmd:metadataStandardName>\r\n        <gco:CharacterString>ISO 19115-2 Geographic information - Metadata - Part 2: Extensions for imagery and gridded data</gco:CharacterString>\r\n      </gmd:metadataStandardName>\r\n      <gmd:metadataStandardVersion>\r\n        <gco:CharacterString>ISO 19115-2:2009(E)</gco:CharacterString>\r\n      </gmd:metadataStandardVersion>\r\n      <gmd:identificationInfo>\r\n        <gmd:MD_DataIdentification>\r\n          <gmd:citation>\r\n            <gmd:CI_Citation>\r\n              <!-- ECS extracts the LongName from here -->\r\n              <!-- UMM-C expects the ShortName to precede the LongName separated by a &gt; here -->\r\n              <gmd:title>\r\n                <gco:CharacterString>ATLAS/ICESat-2 L3A Land and Vegetation Height</gco:CharacterString>\r\n              </gmd:title>\r\n              <gmd:date>\r\n                <gmd:CI_Date>\r\n                  <!-- ECS extracts the RevisionDate from here -->\r\n                  <gmd:date>\r\n                    <gco:Date>2016-06-09</gco:Date>\r\n                  </gmd:date>\r\n                  <gmd:dateType>\r\n                    <gmd:CI_DateTypeCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode\" codeListValue=\"revision\">revision</gmd:CI_DateTypeCode>\r\n                  </gmd:dateType>\r\n                </gmd:CI_Date>\r\n              </gmd:date>\r\n              <!-- VersionID is expected to be here by the Base Reference Metadata Model document -->\r\n              <gmd:edition>\r\n                <gco:CharacterString>003</gco:CharacterString>\r\n              </gmd:edition>\r\n              <gmd:identifier>\r\n                <gmd:MD_Identifier>\r\n                  <!-- ECS extracts the ShortName from here -->\r\n                  <gmd:code>\r\n                    <gco:CharacterString>ATL08</gco:CharacterString>\r\n                  </gmd:code>\r\n                  <gmd:description>\r\n                    <gco:CharacterString>The ECS Short Name</gco:CharacterString>\r\n                  </gmd:description>\r\n                </gmd:MD_Identifier>\r\n              </gmd:identifier>\r\n              <gmd:identifier>\r\n                <gmd:MD_Identifier>\r\n                  <!-- ECS extracts the VersionID from here -->\r\n                  <gmd:code>\r\n                    <gco:CharacterString>003</gco:CharacterString>\r\n                  </gmd:code>\r\n                  <gmd:description>\r\n                    <gco:CharacterString>The ECS Version ID</gco:CharacterString>\r\n                  </gmd:description>\r\n                </gmd:MD_Identifier>\r\n              </gmd:identifier>\r\n              <gmd:identifier>\r\n                <gmd:MD_Identifier>\r\n                  <!-- This field provides the Digital Object Identifier (DOI). -->\r\n                  <gmd:code>\r\n                    <gmx:Anchor xlink:actuate=\"onRequest\" xlink:href=\"http://dx.doi.org/10.5067/ATLAS/ATL08.003\">doi:10.5067/ATLAS/ATL08.003</gmx:Anchor>\r\n                  </gmd:code>\r\n                  <gmd:codeSpace>\r\n                    <gco:CharacterString>gov.nasa.esdis</gco:CharacterString>\r\n                  </gmd:codeSpace>\r\n                  <gmd:description>\r\n                    <gco:CharacterString>A Digital Object Identifier (DOI)</gco:CharacterString>\r\n                  </gmd:description>\r\n                </gmd:MD_Identifier>\r\n              </gmd:identifier>\r\n              <gmd:citedResponsibleParty>\r\n                <gmd:CI_ResponsibleParty>\r\n                  <gmd:organisationName>\r\n                    <gco:CharacterString>National Aeronautics and Space Administration (NASA)</gco:CharacterString>\r\n                  </gmd:organisationName>\r\n                  <gmd:role>\r\n                    <gmd:CI_RoleCode codeList=\"http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_RoleCode\" codeListValue=\"resourceProvider\">resourceProvider</gmd:CI_RoleCode>\r\n                  </gmd:role>\r\n                </gmd:CI_ResponsibleParty>\r\n              </gmd:citedResponsibleParty>\r\n              <gmd:citedResponsibleParty>\r\n                <gmd:CI_ResponsibleParty>\r\n                  <!-- ECS expects ProcessingCenter to be here -->\r\n                  <gmd:organisationName>\r\n                    <gco:CharacterString>GSFC I-SIPS &gt; ICESat-2 Science Investigator-led Processing System</gco:CharacterString>\r\n                  </gmd:organisationName>\r\n                  <gmd:role>\r\n                    <gmd:CI_RoleCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#CI_RoleCode\" codeListValue=\"originator\">originator</gmd:CI_RoleCode>\r\n                  </gmd:role>\r\n                </gmd:CI_ResponsibleParty>\r\n              </gmd:citedResponsibleParty>\r\n              <!-- ECS extracts the VersionDescription from here -->\r\n              <gmd:otherCitationDetails>\r\n                <gco:CharacterString>Initial version of the processing software</gco:CharacterString>\r\n              </gmd:otherCitationDetails>\r\n            </gmd:CI_Citation>\r\n          </gmd:citation>\r\n          <!-- ECS extracts the CollectionDescription from here -->\r\n          <gmd:abstract>\r\n            <gco:CharacterString>The ICESat-2 ATL08 standard data product contains along-track heights of ground and canopy surface at varying length scales. Where data permits, this includes estimates of canopy height, relative canopy cover, canopy height distributions, surface roughness, surface slope/aspect, and apparent reflectance.</gco:CharacterString>\r\n          </gmd:abstract>\r\n          <gmd:purpose>\r\n            <gco:CharacterString>The purpose of ATL08 is to provide along-track land/canopy heights and associated statistics.</gco:CharacterString>\r\n          </gmd:purpose>\r\n          <gmd:credit>\r\n            <gco:CharacterString>The software that generates the ATL08 product was designed and implemented within the ICESat-2 Science Investigator-led Processing System at the NASA Goddard Space Flight Center in Greenbelt, Maryland.</gco:CharacterString>\r\n          </gmd:credit>\r\n          <gmd:status>\r\n            <gmd:MD_ProgressCode codeList=\"http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_ProgressCode\" codeListValue=\"onGoing\">onGoing</gmd:MD_ProgressCode>\r\n          </gmd:status>\r\n          <gmd:pointOfContact>\r\n            <gmd:CI_ResponsibleParty>\r\n              <!-- ECS expects ArchiveCenter to be here -->\r\n              <gmd:organisationName>\r\n                <gco:CharacterString>NSIDC DAAC &gt; NASA National Snow and Ice Data Center Distributed Active Archive Center</gco:CharacterString>\r\n              </gmd:organisationName>\r\n              <gmd:contactInfo xlink:href=\"#NSIDC_DAAC_CONTACT_ID\"/>\r\n              <gmd:role>\r\n                <gmd:CI_RoleCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#CI_RoleCode\" codeListValue=\"distributor\">distributor</gmd:CI_RoleCode>\r\n              </gmd:role>\r\n            </gmd:CI_ResponsibleParty>\r\n          </gmd:pointOfContact>\r\n          <gmd:resourceFormat>\r\n            <gmd:MD_Format>\r\n              <gmd:name>\r\n                <gco:CharacterString>HDF</gco:CharacterString>\r\n              </gmd:name>\r\n              <gmd:version>\r\n                <gco:CharacterString>5</gco:CharacterString>\r\n              </gmd:version>\r\n            </gmd:MD_Format>\r\n          </gmd:resourceFormat>\r\n          <gmd:descriptiveKeywords>\r\n            <gmd:MD_Keywords>\r\n              <gmd:keyword>\r\n                <gco:CharacterString>EARTH SCIENCE &gt; BIOSPHERE &gt; VEGETATION &gt; NONE &gt; NONE &gt; NONE &gt; NONE</gco:CharacterString>\r\n              </gmd:keyword>\r\n              <gmd:keyword>\r\n                <gco:CharacterString>EARTH SCIENCE &gt; BIOSPHERE &gt; VEGETATION &gt; VEGETATION COVER &gt; NONE &gt; NONE &gt; NONE</gco:CharacterString>\r\n              </gmd:keyword>\r\n              <gmd:keyword>\r\n                <gco:CharacterString>EARTH SCIENCE &gt; LAND SURFACE &gt; NONE &gt; NONE &gt; NONE &gt; NONE &gt; NONE</gco:CharacterString>\r\n              </gmd:keyword>\r\n              <gmd:keyword>\r\n                <gco:CharacterString>EARTH SCIENCE &gt; LAND SURFACE &gt; TOPOGRAPHY &gt; SURFACE ROUGHNESS &gt; NONE &gt; NONE &gt; NONE</gco:CharacterString>\r\n              </gmd:keyword>\r\n              <gmd:keyword>\r\n                <gco:CharacterString>EARTH SCIENCE &gt; LAND SURFACE &gt; TOPOGRAPHY &gt; TERRAIN ELEVATION &gt; NONE &gt; NONE &gt; NONE</gco:CharacterString>\r\n              </gmd:keyword>\r\n              <gmd:type>\r\n                <gmd:MD_KeywordTypeCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#MD_KeywordTypeCode\" codeListValue=\"theme\">theme</gmd:MD_KeywordTypeCode>\r\n              </gmd:type>\r\n              <gmd:thesaurusName>\r\n                <gmd:CI_Citation>\r\n                  <gmd:title>\r\n                    <gco:CharacterString>NASA/GCMD Science Keywords</gco:CharacterString>\r\n                  </gmd:title>\r\n                  <gmd:date gco:nilReason=\"unknown\"/>\r\n                  <gmd:citedResponsibleParty>\r\n                    <gmd:CI_ResponsibleParty id=\"GCMD_USO_ID\">\r\n                      <gmd:organisationName>\r\n                        <gco:CharacterString>NASA Global Change Master Directory (GCMD) User Support Office</gco:CharacterString>\r\n                      </gmd:organisationName>\r\n                      <gmd:contactInfo>\r\n                        <gmd:CI_Contact>\r\n                          <gmd:phone gco:nilReason=\"missing\"/>\r\n                          <gmd:address>\r\n                            <gmd:CI_Address>\r\n                              <gmd:deliveryPoint>\r\n                                <gco:CharacterString>NASA Global Change Master Directory, Goddard Space Flight Center</gco:CharacterString>\r\n                              </gmd:deliveryPoint>\r\n                              <gmd:city>\r\n                                <gco:CharacterString>Greenbelt</gco:CharacterString>\r\n                              </gmd:city>\r\n                              <gmd:administrativeArea>\r\n                                <gco:CharacterString>MD</gco:CharacterString>\r\n                              </gmd:administrativeArea>\r\n                              <gmd:postalCode>\r\n                                <gco:CharacterString>20771</gco:CharacterString>\r\n                              </gmd:postalCode>\r\n                              <gmd:country>\r\n                                <gco:CharacterString>USA</gco:CharacterString>\r\n                              </gmd:country>\r\n                              <gmd:electronicMailAddress>\r\n                                <gco:CharacterString>gcmduso@gcmd.gsfc.nasa.gov</gco:CharacterString>\r\n                              </gmd:electronicMailAddress>\r\n                            </gmd:CI_Address>\r\n                          </gmd:address>\r\n                          <gmd:onlineResource>\r\n                            <gmd:CI_OnlineResource>\r\n                              <gmd:linkage>\r\n                                <gmd:URL>http://gcmd.nasa.gov/</gmd:URL>\r\n                              </gmd:linkage>\r\n                              <gmd:protocol>\r\n                                <gco:CharacterString>http</gco:CharacterString>\r\n                              </gmd:protocol>\r\n                              <gmd:applicationProfile>\r\n                                <gco:CharacterString>web browser</gco:CharacterString>\r\n                              </gmd:applicationProfile>\r\n                              <gmd:name>\r\n                                <gco:CharacterString>NASA Global Change Master Directory (GCMD)</gco:CharacterString>\r\n                              </gmd:name>\r\n                              <gmd:description>\r\n                                <gco:CharacterString>Home Page</gco:CharacterString>\r\n                              </gmd:description>\r\n                              <gmd:function>\r\n                                <gmd:CI_OnLineFunctionCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#CI_OnLineFunctionCode\" codeListValue=\"information\">information</gmd:CI_OnLineFunctionCode>\r\n                              </gmd:function>\r\n                            </gmd:CI_OnlineResource>\r\n                          </gmd:onlineResource>\r\n                          <gmd:contactInstructions>\r\n                            <gco:CharacterString>http://gcmd.nasa.gov/MailComments/MailComments.jsf?rcpt=gcmduso</gco:CharacterString>\r\n                          </gmd:contactInstructions>\r\n                        </gmd:CI_Contact>\r\n                      </gmd:contactInfo>\r\n                      <gmd:role>\r\n                        <gmd:CI_RoleCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#CI_RoleCode\" codeListValue=\"custodian\">custodian</gmd:CI_RoleCode>\r\n                      </gmd:role>\r\n                    </gmd:CI_ResponsibleParty>\r\n                  </gmd:citedResponsibleParty>\r\n                  <gmd:citedResponsibleParty>\r\n                    <gmd:CI_ResponsibleParty id=\"GCMD_KEYWORDS_ID\">\r\n                      <gmd:organisationName>\r\n                        <gco:CharacterString>Global Change Master Directory (GCMD)</gco:CharacterString>\r\n                      </gmd:organisationName>\r\n                      <gmd:contactInfo>\r\n                        <gmd:CI_Contact>\r\n                          <gmd:phone gco:nilReason=\"missing\"/>\r\n                          <gmd:address>\r\n                            <gmd:CI_Address>\r\n                              <gmd:deliveryPoint>\r\n                                <gco:CharacterString>NASA Global Change Master Directory, Goddard Space Flight Center</gco:CharacterString>\r\n                              </gmd:deliveryPoint>\r\n                              <gmd:city>\r\n                                <gco:CharacterString>Greenbelt</gco:CharacterString>\r\n                              </gmd:city>\r\n                              <gmd:administrativeArea>\r\n                                <gco:CharacterString>MD</gco:CharacterString>\r\n                              </gmd:administrativeArea>\r\n                              <gmd:postalCode>\r\n                                <gco:CharacterString>20771</gco:CharacterString>\r\n                              </gmd:postalCode>\r\n                              <gmd:country>\r\n                                <gco:CharacterString>USA</gco:CharacterString>\r\n                              </gmd:country>\r\n                              <gmd:electronicMailAddress>\r\n                                <gco:CharacterString>gcmduso@gcmd.gsfc.nasa.gov</gco:CharacterString>\r\n                              </gmd:electronicMailAddress>\r\n                            </gmd:CI_Address>\r\n                          </gmd:address>\r\n                          <gmd:onlineResource>\r\n                            <gmd:CI_OnlineResource>\r\n                              <gmd:linkage>\r\n                                <gmd:URL>http://gcmd.nasa.gov/Resources/valids/</gmd:URL>\r\n                              </gmd:linkage>\r\n                              <gmd:protocol>\r\n                                <gco:CharacterString>http</gco:CharacterString>\r\n                              </gmd:protocol>\r\n                              <gmd:applicationProfile>\r\n                                <gco:CharacterString>web browser</gco:CharacterString>\r\n                              </gmd:applicationProfile>\r\n                              <gmd:name>\r\n                                <gco:CharacterString>NASA Global Change Master Directory (GCMD) Keyword Page</gco:CharacterString>\r\n                              </gmd:name>\r\n                              <gmd:description>\r\n                                <gco:CharacterString>This page describes the NASA GCMD Keywords, how to reference those keywords and provides download instructions.</gco:CharacterString>\r\n                              </gmd:description>\r\n                              <gmd:function>\r\n                                <gmd:CI_OnLineFunctionCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#CI_OnLineFunctionCode\" codeListValue=\"download\">download</gmd:CI_OnLineFunctionCode>\r\n                              </gmd:function>\r\n                            </gmd:CI_OnlineResource>\r\n                          </gmd:onlineResource>\r\n                          <gmd:contactInstructions>\r\n                            <gco:CharacterString>http://gcmd.nasa.gov/MailComments/MailComments.jsf?rcpt=gcmduso</gco:CharacterString>\r\n                          </gmd:contactInstructions>\r\n                        </gmd:CI_Contact>\r\n                      </gmd:contactInfo>\r\n                      <gmd:role>\r\n                        <gmd:CI_RoleCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#CI_RoleCode\" codeListValue=\"custodian\">custodian</gmd:CI_RoleCode>\r\n                      </gmd:role>\r\n                    </gmd:CI_ResponsibleParty>\r\n                  </gmd:citedResponsibleParty>\r\n                </gmd:CI_Citation>\r\n              </gmd:thesaurusName>\r\n            </gmd:MD_Keywords>\r\n          </gmd:descriptiveKeywords>\r\n          <gmd:descriptiveKeywords>\r\n            <gmd:MD_Keywords>\r\n              <gmd:keyword>\r\n                <gco:CharacterString>GEOGRAPHIC REGION &gt; GLOBAL</gco:CharacterString>\r\n              </gmd:keyword>\r\n              <gmd:type>\r\n                <gmd:MD_KeywordTypeCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#MD_KeywordTypeCode\" codeListValue=\"place\">place</gmd:MD_KeywordTypeCode>\r\n              </gmd:type>\r\n              <gmd:thesaurusName>\r\n                <gmd:CI_Citation>\r\n                  <gmd:title>\r\n                    <gco:CharacterString>NASA/GCMD Location Keywords</gco:CharacterString>\r\n                  </gmd:title>\r\n                  <gmd:date gco:nilReason=\"unknown\"/>\r\n                  <gmd:citedResponsibleParty xlink:href=\"#GCMD_USO_ID\"/>\r\n                  <gmd:citedResponsibleParty xlink:href=\"#GCMD_KEYWORDS_ID\"/>\r\n                </gmd:CI_Citation>\r\n              </gmd:thesaurusName>\r\n            </gmd:MD_Keywords>\r\n          </gmd:descriptiveKeywords>\r\n          <gmd:descriptiveKeywords>\r\n            <gmd:MD_Keywords>\r\n              <gmd:keyword>\r\n                <gco:CharacterString>NASA/NSIDC_DAAC &gt; NASA National Snow and Ice Data Center Distributed Active Archive Center</gco:CharacterString>\r\n              </gmd:keyword>\r\n              <gmd:type>\r\n                <gmd:MD_KeywordTypeCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#MD_KeywordTypeCode\" codeListValue=\"dataCenter\">dataCenter</gmd:MD_KeywordTypeCode>\r\n              </gmd:type>\r\n              <gmd:thesaurusName>\r\n                <gmd:CI_Citation>\r\n                  <gmd:title>\r\n                    <gco:CharacterString>NASA/GCMD Data Center Keywords</gco:CharacterString>\r\n                  </gmd:title>\r\n                  <gmd:date gco:nilReason=\"unknown\"/>\r\n                  <gmd:citedResponsibleParty xlink:href=\"#GCMD_USO_ID\"/>\r\n                  <gmd:citedResponsibleParty xlink:href=\"#GCMD_KEYWORDS_ID\"/>\r\n                </gmd:CI_Citation>\r\n              </gmd:thesaurusName>\r\n            </gmd:MD_Keywords>\r\n          </gmd:descriptiveKeywords>\r\n          <gmd:descriptiveKeywords>\r\n            <gmd:MD_Keywords>\r\n              <gmd:keyword>\r\n                <gco:CharacterString>Earth Observation Satellites &gt; NASA Decadal Survey &gt; ICESAT-2 &gt; Ice, Cloud, and land Elevation Satellite-2</gco:CharacterString>\r\n              </gmd:keyword>\r\n              <gmd:type>\r\n                <gmd:MD_KeywordTypeCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#MD_KeywordTypeCode\" codeListValue=\"platform\">platform</gmd:MD_KeywordTypeCode>\r\n              </gmd:type>\r\n              <gmd:thesaurusName>\r\n                <gmd:CI_Citation>\r\n                  <gmd:title>\r\n                    <gco:CharacterString>NASA/GCMD Platform Keywords</gco:CharacterString>\r\n                  </gmd:title>\r\n                  <gmd:date gco:nilReason=\"unknown\"/>\r\n                  <gmd:citedResponsibleParty xlink:href=\"#GCMD_USO_ID\"/>\r\n                  <gmd:citedResponsibleParty xlink:href=\"#GCMD_KEYWORDS_ID\"/>\r\n                </gmd:CI_Citation>\r\n              </gmd:thesaurusName>\r\n            </gmd:MD_Keywords>\r\n          </gmd:descriptiveKeywords>\r\n          <gmd:descriptiveKeywords>\r\n            <gmd:MD_Keywords>\r\n              <gmd:keyword>\r\n                <gco:CharacterString>Earth Remote Sensing Instruments &gt; Active Remote Sensing &gt; Altimeters &gt; Lidar/Laser Altimeters &gt; ATLAS &gt; Advanced Topographic Laser Altimeter System</gco:CharacterString>\r\n              </gmd:keyword>\r\n              <gmd:type>\r\n                <gmd:MD_KeywordTypeCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#MD_KeywordTypeCode\" codeListValue=\"instrument\">instrument</gmd:MD_KeywordTypeCode>\r\n              </gmd:type>\r\n              <gmd:thesaurusName>\r\n                <gmd:CI_Citation>\r\n                  <gmd:title>\r\n                    <gco:CharacterString>NASA/GCMD Instrument Keywords</gco:CharacterString>\r\n                  </gmd:title>\r\n                  <gmd:date gco:nilReason=\"unknown\"/>\r\n                  <gmd:citedResponsibleParty xlink:href=\"#GCMD_USO_ID\"/>\r\n                  <gmd:citedResponsibleParty xlink:href=\"#GCMD_KEYWORDS_ID\"/>\r\n                </gmd:CI_Citation>\r\n              </gmd:thesaurusName>\r\n            </gmd:MD_Keywords>\r\n          </gmd:descriptiveKeywords>\r\n          <gmd:resourceConstraints>\r\n            <gmd:MD_Constraints>\r\n              <gmd:useLimitation>\r\n                <gco:CharacterString>Cite these data in publications as follows: The data used in this study were produced by the ICESat-2 Science Project Office at NASA/GSFC. The data archive site is the NASA National Snow and Ice Data Center Distributed Active Archive Center.</gco:CharacterString>\r\n              </gmd:useLimitation>\r\n            </gmd:MD_Constraints>\r\n          </gmd:resourceConstraints>\r\n          <gmd:language>\r\n            <gco:CharacterString>eng</gco:CharacterString>\r\n          </gmd:language>\r\n          <gmd:topicCategory>\r\n            <gmd:MD_TopicCategoryCode>geoscientificInformation</gmd:MD_TopicCategoryCode>\r\n          </gmd:topicCategory>\r\ni          <gmd:extent>\r\n            <gmd:EX_Extent id=\"boundingExtent\">\r\n              <gmd:description>\r\n                <gco:CharacterString>SpatialCoverageType=HORIZONTAL, SpatialGranuleSpatialRepresentation=ORBIT, TemporalRangeType=Continuous Range, TimeType=UTC</gco:CharacterString>\r\n              </gmd:description>\r\n              <gmd:geographicElement>\r\n                <gmd:EX_GeographicBoundingBox>\r\n                  <!-- ECS extracts WestBoundingCoordinate from here -->\r\n                  <gmd:westBoundLongitude>\r\n                    <gco:Decimal>-180.0</gco:Decimal>\r\n                  </gmd:westBoundLongitude>\r\n                  <!-- ECS extracts EastBoundingCoordinate from here -->\r\n                  <gmd:eastBoundLongitude>\r\n                    <gco:Decimal>180.0</gco:Decimal>\r\n                  </gmd:eastBoundLongitude>\r\n                  <!-- ECS extracts SouthBoundingCoordinate from here -->\r\n                  <gmd:southBoundLatitude>\r\n                    <gco:Decimal>-90.0</gco:Decimal>\r\n                  </gmd:southBoundLatitude>\r\n                  <!-- ECS extracts NorthBoundingCoordinate from here -->\r\n                  <gmd:northBoundLatitude>\r\n                    <gco:Decimal>90.0</gco:Decimal>\r\n                  </gmd:northBoundLatitude>\r\n                </gmd:EX_GeographicBoundingBox>\r\n              </gmd:geographicElement>\r\n              <gmd:geographicElement>\r\n                <gmd:EX_GeographicDescription>\r\n                  <gmd:geographicIdentifier>\r\n                    <gmd:MD_Identifier>\r\n                      <gmd:code>\r\n                        <gco:CharacterString>SwathWidth: 36.0 Period: 96.8 InclinationAngle: 92.0 NumberOfOrbits: 0.071428571 StartCircularLatitude: 0.0</gco:CharacterString>\r\n                      </gmd:code>\r\n                      <gmd:codeSpace>\r\n                        <gco:CharacterString>gov.nasa.esdis.umm.orbitparameters</gco:CharacterString>\r\n                      </gmd:codeSpace>\r\n                      <gmd:description>\r\n                        <gco:CharacterString>OrbitParameters</gco:CharacterString>\r\n                      </gmd:description>\r\n                    </gmd:MD_Identifier>\r\n                  </gmd:geographicIdentifier>\r\n                </gmd:EX_GeographicDescription>\r\n              </gmd:geographicElement>\r\n              <gmd:temporalElement>\r\n                <gmd:EX_TemporalExtent>\r\n                  <gmd:extent>\r\n                    <gml:TimePeriod gml:id=\"TimePeriod_ID_1\">\r\n                      <!-- ECS extracts RangeBeginningDate and RangeBeginningTime from here -->\r\n                      <gml:beginPosition>2005-01-01T00:00:00Z</gml:beginPosition>\r\n                      <!-- ECS extracts RangeEndingDate and RangeEndingTime from here -->\r\n                      <gml:endPosition>2020-12-31T23:59:59Z</gml:endPosition>\r\n                    </gml:TimePeriod>\r\n                  </gmd:extent>\r\n                </gmd:EX_TemporalExtent>\r\n              </gmd:temporalElement>\r\n            </gmd:EX_Extent>\r\n          </gmd:extent>\r\n          <gmd:processingLevel>\r\n            <gmd:MD_Identifier>\r\n              <gmd:code>\r\n                <gco:CharacterString>3A</gco:CharacterString>\r\n              </gmd:code>\r\n              <gmd:description gco:nilReason=\"missing\"/>\r\n            </gmd:MD_Identifier>\r\n          </gmd:processingLevel>\r\n        </gmd:MD_DataIdentification>\r\n      </gmd:identificationInfo>\r\n      <gmd:contentInfo>\r\n        <gmd:MD_ImageDescription>\r\n          <gmd:attributeDescription gco:nilReason=\"missing\"/>\r\n          <gmd:contentType gco:nilReason=\"missing\"/>\r\n          <gmd:processingLevelCode>\r\n            <gmd:MD_Identifier>\r\n              <gmd:code>\r\n                <gco:CharacterString>3A</gco:CharacterString>\r\n              </gmd:code>\r\n              <gmd:description gco:nilReason=\"missing\"/>\r\n            </gmd:MD_Identifier>\r\n          </gmd:processingLevelCode>\r\n        </gmd:MD_ImageDescription>\r\n      </gmd:contentInfo>\r\n      <gmd:distributionInfo>\r\n        <gmd:MD_Distribution>\r\n          <gmd:distributionFormat>\r\n            <gmd:MD_Format>\r\n              <gmd:name>\r\n                <gco:CharacterString>HDF</gco:CharacterString>\r\n              </gmd:name>\r\n              <gmd:version>\r\n                <gco:CharacterString>5</gco:CharacterString>\r\n              </gmd:version>\r\n            </gmd:MD_Format>\r\n          </gmd:distributionFormat>\r\n          <gmd:distributor>\r\n            <gmd:MD_Distributor>\r\n              <gmd:distributorContact>\r\n                <gmd:CI_ResponsibleParty>\r\n                  <gmd:organisationName>\r\n                    <gco:CharacterString>NSIDC DAAC &gt; NASA National Snow and Ice Data Center Distributed Active Archive Center</gco:CharacterString>\r\n                  </gmd:organisationName>\r\n                  <gmd:contactInfo xlink:href=\"#NSIDC_DAAC_CONTACT_ID\"/>\r\n                  <gmd:role>\r\n                    <gmd:CI_RoleCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#CI_RoleCode\" codeListValue=\"distributor\">distributor</gmd:CI_RoleCode>\r\n                  </gmd:role>\r\n                </gmd:CI_ResponsibleParty>\r\n              </gmd:distributorContact>\r\n              <gmd:distributorTransferOptions>\r\n                <gmd:MD_DigitalTransferOptions>\r\n                  <gmd:onLine>\r\n                    <gmd:CI_OnlineResource>\r\n                      <gmd:linkage>\r\n                        <gmd:URL>http://nsidc.org/data/icesat2/data.html</gmd:URL>\r\n                      </gmd:linkage>\r\n                      <gmd:protocol>\r\n                        <gco:CharacterString>http</gco:CharacterString>\r\n                      </gmd:protocol>\r\n                      <gmd:description>\r\n                        <gco:CharacterString>Data Product Description Page</gco:CharacterString>\r\n                      </gmd:description>\r\n                      <gmd:function>\r\n                        <gmd:CI_OnLineFunctionCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#CI_OnLineFunctionCode\" codeListValue=\"information\">information</gmd:CI_OnLineFunctionCode>\r\n                      </gmd:function>\r\n                    </gmd:CI_OnlineResource>\r\n                  </gmd:onLine>\r\n                  <gmd:onLine>\r\n                    <gmd:CI_OnlineResource>\r\n                      <gmd:linkage>\r\n                        <gmd:URL>http://nsidc.org/data/icesat2/order.html</gmd:URL>\r\n                      </gmd:linkage>\r\n                      <gmd:protocol>\r\n                        <gco:CharacterString>http</gco:CharacterString>\r\n                      </gmd:protocol>\r\n                      <gmd:description>\r\n                        <gco:CharacterString>Data Product Order Page</gco:CharacterString>\r\n                      </gmd:description>\r\n                      <gmd:function>\r\n                        <gmd:CI_OnLineFunctionCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#CI_OnLineFunctionCode\" codeListValue=\"order\">order</gmd:CI_OnLineFunctionCode>\r\n                      </gmd:function>\r\n                    </gmd:CI_OnlineResource>\r\n                  </gmd:onLine>\r\n                  <gmd:onLine>\r\n                    <gmd:CI_OnlineResource>\r\n                      <gmd:linkage>\r\n                        <gmd:URL>http://dx.doi.org/10.5067/ATLAS/ATL08.003</gmd:URL>\r\n                      </gmd:linkage>\r\n                      <gmd:protocol>\r\n                        <gco:CharacterString>http</gco:CharacterString>\r\n                      </gmd:protocol>\r\n                      <gmd:description>\r\n                        <gco:CharacterString>Digital Object Identifier URL</gco:CharacterString>\r\n                      </gmd:description>\r\n                      <gmd:function>\r\n                        <gmd:CI_OnLineFunctionCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#CI_OnLineFunctionCode\" codeListValue=\"information\">information</gmd:CI_OnLineFunctionCode>\r\n                      </gmd:function>\r\n                    </gmd:CI_OnlineResource>\r\n                  </gmd:onLine>\r\n                </gmd:MD_DigitalTransferOptions>\r\n              </gmd:distributorTransferOptions>\r\n            </gmd:MD_Distributor>\r\n          </gmd:distributor>\r\n        </gmd:MD_Distribution>\r\n      </gmd:distributionInfo>\r\n      <gmi:acquisitionInformation>\r\n        <gmi:MI_AcquisitionInformation>\r\n          <gmi:instrument>\r\n            <eos:EOS_Instrument id=\"ATLAS_INSTRUMENT_ID\">\r\n              <gmi:citation>\r\n                <gmd:CI_Citation>\r\n                  <gmd:title>\r\n                    <gco:CharacterString>ATLAS &gt; Advanced Topographic Laser Altimeter System</gco:CharacterString>\r\n                  </gmd:title>\r\n                  <gmd:date gco:nilReason=\"unknown\"/>\r\n                </gmd:CI_Citation>\r\n              </gmi:citation>\r\n              <gmi:identifier>\r\n                <gmd:MD_Identifier>\r\n                  <gmd:code>\r\n                    <gco:CharacterString>ATLAS</gco:CharacterString>\r\n                  </gmd:code>\r\n                  <gmd:description>\r\n                    <gco:CharacterString>Advanced Topographic Laser Altimeter System</gco:CharacterString>\r\n                  </gmd:description>\r\n                </gmd:MD_Identifier>\r\n              </gmi:identifier>\r\n              <gmi:type>\r\n                <gco:CharacterString>Laser Altimeter</gco:CharacterString>\r\n              </gmi:type>\r\n              <gmi:description>\r\n                <gco:CharacterString>ATLAS on ICESat-2 determines the range between the satellite and the Earth\'s surface by measuring the two-way time delay of short pulses of laser light that it transmits in six beams.  It is different from previous operational ice-sheet altimeters in that it is a photon-counting LIDAR.  ATLAS records a set of arrival times for individual photons, which are then analyzed to derive surface, vegetation, and cloud properties.  ATLAS has six beams arranged in three pairs, so that it samples each of three reference pair tracks with a pair of beams; ATLAS transmits pulses at 10 kHz, giving approximately one pulse every 0.7 m along track; ATLAS\'s expected pointing control will be better than 90 m RMS.</gco:CharacterString>\r\n              </gmi:description>\r\n              <gmi:mountedOn xlink:href=\"#ICESAT_2_PLATFORM_ID\"/>\r\n            </eos:EOS_Instrument>\r\n          </gmi:instrument>\r\n          <gmi:operation>\r\n            <!-- MI_Operation is expected to be here by the Base Reference Metadata Model document-->\r\n            <gmi:MI_Operation>\r\n              <gmi:description>\r\n                <gco:CharacterString>ICESat-2 &gt; Ice, Cloud, and land Elevation Satellite-2</gco:CharacterString>\r\n              </gmi:description>\r\n              <gmi:citation>\r\n                <gmd:CI_Citation>\r\n                  <gmd:title>\r\n                    <gco:CharacterString>ICESat-2 &gt; Ice, Cloud, and land Elevation Satellite-2</gco:CharacterString>\r\n                  </gmd:title>\r\n                  <gmd:date gco:nilReason=\"unknown\"/>\r\n                </gmd:CI_Citation>\r\n              </gmi:citation>\r\n              <gmi:identifier>\r\n                <gmd:MD_Identifier>\r\n                  <gmd:code>\r\n                    <gco:CharacterString>ICESat-2</gco:CharacterString>\r\n                  </gmd:code>\r\n                  <gmd:description>\r\n                    <gco:CharacterString>Ice, Cloud, and land Elevation Satellite-2</gco:CharacterString>\r\n                  </gmd:description>\r\n                </gmd:MD_Identifier>\r\n              </gmi:identifier>\r\n              <gmi:status>\r\n                <gmd:MD_ProgressCode codeList=\"http://cdn.earthdata.nasa.gov/iso/resources/Codelist/gmxCodelists.xml#MD_ProgressCode\" codeListValue=\"underDevelopment\">underDevelopment</gmd:MD_ProgressCode>\r\n              </gmi:status>\r\n              <gmi:parentOperation gco:nilReason=\"inapplicable\"/>\r\n              <gmi:platform xlink:href=\"#ICESAT_2_PLATFORM_ID\"/>\r\n            </gmi:MI_Operation>\r\n          </gmi:operation>\r\n          <gmi:platform>\r\n            <eos:EOS_Platform id=\"ICESAT_2_PLATFORM_ID\">\r\n              <gmi:citation>\r\n                <gmd:CI_Citation>\r\n                  <gmd:title>\r\n                    <gco:CharacterString>ICESat-2 &gt; Ice, Cloud, and land Elevation Satellite-2</gco:CharacterString>\r\n                  </gmd:title>\r\n                  <gmd:date gco:nilReason=\"unknown\"/>\r\n                </gmd:CI_Citation>\r\n              </gmi:citation>\r\n              <gmi:identifier>\r\n                <gmd:MD_Identifier>\r\n                  <gmd:code>\r\n                    <gco:CharacterString>ICESat-2</gco:CharacterString>\r\n                  </gmd:code>\r\n                  <gmd:description>\r\n                    <gco:CharacterString>Ice, Cloud, and land Elevation Satellite-2</gco:CharacterString>\r\n                  </gmd:description>\r\n                </gmd:MD_Identifier>\r\n              </gmi:identifier>\r\n              <gmi:description>\r\n                <gco:CharacterString>Spacecraft</gco:CharacterString>\r\n              </gmi:description>\r\n              <gmi:instrument xlink:href=\"#ATLAS_INSTRUMENT_ID\"/>\r\n            </eos:EOS_Platform>\r\n          </gmi:platform>\r\n        </gmi:MI_AcquisitionInformation>\r\n      </gmi:acquisitionInformation>\r\n    </gmi:MI_Metadata>\r\n  </gmd:seriesMetadata>\r\n</gmd:DS_Series>\r\n" ;

  group: AcquisitionInformation {

    group: lidar {

      // group attributes:
      		:pulse_rate = "10000 pps" ;
      		:wavelength = "532 nm" ;
      		:identifier = "ATLAS" ;
      		:type = "Laser Altimeter" ;
      		:description = "ATLAS on ICESat-2 determines the range between the satellite and the Earth\'s surface by measuring the two-way time delay of short pulses of laser light that it transmits in six beams.  It is different from previous operational ice-sheet altimeters in that it is a photon-counting LIDAR.  ATLAS records a set of arrival times for individual photons, which are then analyzed to derive surface, vegetation, and cloud properties.  ATLAS has six beams arranged in three pairs, so that it samples each of three reference pair tracks with a pair of beams; ATLAS transmits pulses at 10 kHz, giving approximately one pulse every 0.7 m along track; ATLAS\'s expected pointing control will be better than 90 m RMS." ;
      } // group lidar

    group: lidarDocument {

      // group attributes:
      		:edition = "Pre-Release" ;
      		:publicationDate = "12/31/17" ;
      		:title = "A document describing the ATLAS instrument will be provided by the ICESat-2 Project Science Office." ;
      } // group lidarDocument

    group: platform {

      // group attributes:
      		:identifier = "ICESat-2" ;
      		:description = "Ice, Cloud, and land Elevation Satellite-2" ;
      		:type = "Spacecraft" ;
      } // group platform

    group: platformDocument {

      // group attributes:
      		:edition = "31-Dec-16" ;
      		:publicationDate = "31-Dec-16" ;
      		:title = "The Ice, Cloud, and land Elevation Satellite-2 (ICESat-2): Science requirements, concept, and implementation. Thorsten Markus, Tom Neumann, Anthony Martino, Waleed Abdalati, Kelly Brunt, Beata Csatho, Sinead Farrell, Helen Fricker, Alex Gardner, David Harding, Michael Jasinski, Ron Kwok, Lori Magruder, Dan Lubin, Scott Luthcke, James Morison, Ross Nelson, Amy Neuenschwander, Stephen Palm, Sorin Popescu, CK Shum, Bob E. Schutz, Benjamin Smith, Yuekui Yang, Jay Zwally. http://dx.doi.org/10.1016/j.rse.2016.12.029" ;
      } // group platformDocument
    } // group AcquisitionInformation

  group: DataQuality {

    // group attributes:
    		:scope = "NOT_SET" ;

    group: CompletenessOmission {

      // group attributes:
      		:evaluationMethodType = "directInternal" ;
      		:measureDescription = "TBD" ;
      		:nameOfMeasure = "TBD" ;
      		:unitofMeasure = "TBD" ;
      		:value = "NOT_SET" ;
      } // group CompletenessOmission

    group: DomainConsistency {

      // group attributes:
      		:evaluationMethodType = "directInternal" ;
      		:measureDescription = "TBD" ;
      		:nameOfMeasure = "TBD" ;
      		:unitofMeasure = "TBD" ;
      		:value = "NOT_SET" ;
      } // group DomainConsistency
    } // group DataQuality

  group: DatasetIdentification {

    // group attributes:
    		:spatialRepresentationType = "along-track" ;
    		:creationDate = "2020-04-01T14:03:26.000000Z" ;
    		:uuid = "ae899cbd-cf20-3541-9952-cb5220d5467b" ;
    		:fileName = "ATL08_20181014084920_02400109_003_01.h5" ;
    		:VersionID = "003" ;
    		:language = "eng" ;
    		:characterSet = "utf8" ;
    		:shortName = "ATL08" ;
    		:originatorOrganizationName = "GSFC I-SIPS > ICESat-2 Science Investigator-led Processing System" ;
    		:abstract = "The ICESat-2 ATL08 standard data product contains along-track heights of ground and canopy surface at varying length scales. Where data permits, this includes estimates of canopy height, relative canopy cover, canopy height distributions, surface roughness, surface slope/aspect, and apparent reflectance." ;
    		:purpose = "The purpose of ATL08 is to provide along-track land/canopy heights and associated statistics." ;
    		:credit = "The software that generates the ATL08 product was designed and implemented within the ICESat-2 Science Investigator-led Processing System at the NASA Goddard Space Flight Center in Greenbelt, Maryland." ;
    		:status = "onGoing" ;
    		:topicCategory = "geoscientificInformation" ;
    } // group DatasetIdentification

  group: Extent {

    // group attributes:
    		:northBoundLatitude = -33.6666200966049 ;
    		:eastBoundLongitude = -80.4274386927379 ;
    		:southBoundLatitude = -33.6709309916173 ;
    		:westBoundLongitude = -80.4279359434023 ;
    		:rangeBeginningDateTime = "2018-10-14T08:51:05.104949Z" ;
    		:rangeEndingDateTime = "2018-10-14T08:51:05.172649Z" ;
    } // group Extent

  group: Lineage {

    group: ANC06-01 {

      // group attributes:
      		:description = "GMTED 7.5 arcsec Digital Elevation Model reformatted into HDF5 and re-referenced to the WGS-84 ellipsoid." ;
      		:fileName = "gmted75_20180705_001_01.h5" ;
      		:shortName = "ANC06-01" ;
      		:uuid = "a44debc8-29af-3744-860c-227b37a4da6f" ;
      		:version = "20180705" ;
      } // group ANC06-01

    group: ANC06-02 {

      // group attributes:
      		:description = "ArcticDEM 32m Digital Elevation Model reformatted into HDF5." ;
      		:fileName = "arcticdem32m_20190611_001_01.h5" ;
      		:shortName = "ANC06-02" ;
      		:uuid = "ce07ef72-0bf4-353b-8475-fb568b029905" ;
      		:version = "20190611" ;
      } // group ANC06-02

    group: ANC06-03 {

      // group attributes:
      		:description = "REMA Antarctica 100m Digital Elevation Model filled and reformatted into HDF5" ;
      		:fileName = "atl06rema100m_20190628_001_01.h5" ;
      		:shortName = "ANC06-03" ;
      		:uuid = "3e0a81bd-bbd5-35fa-b868-3254f9355b7f" ;
      		:version = "20190628" ;
      } // group ANC06-03

    group: ANC14 {

      // group attributes:
      		:description = "Landsat Canopy Mask File" ;
      		:fileName = "" ;
      		:shortName = "ANC14" ;
      		:uuid = "" ;
      		:version = "" ;
      } // group ANC14

    group: ANC18 {

      // group attributes:
      		:description = "Modis Land Cover Mask File" ;
      		:fileName = "glcc_2012_20180226_001_global.h5" ;
      		:shortName = "ANC18" ;
      		:uuid = "46e34ac9-892a-3a9d-ab7e-6a329e167a1a" ;
      		:version = "20180226" ;
      } // group ANC18

    group: ANC19 {

      // group attributes:
      		:description = "TAI to UTC leapsecond file retrieved from ftp://maia.usno.navy.mil/ser7/tai-utc.dat" ;
      		:fileName = "tai_utc_2017.dat" ;
      		:shortName = "ANC19" ;
      		:uuid = "7c66d365-278a-31f7-8fe4-9c80e2f012e5" ;
      		:version = "001" ;
      } // group ANC19

    group: ANC25-08 {

      // group attributes:
      		:description = "HDF5 template file that defines the organization and default content of the product." ;
      		:fileName = "ANC25-08_20200311154328_033_01.h5" ;
      		:shortName = "ANC25-08" ;
      		:uuid = "654d3fff-958d-3dbe-8f73-ca718a5538fd" ;
      		:version = "033" ;
      } // group ANC25-08

    group: ANC26-08 {

      // group attributes:
      		:description = "HDF5 template file that defines the organization and default content of the product metadata." ;
      		:fileName = "ANC26-08_20200311154329_033_01.h5" ;
      		:shortName = "ANC26-08" ;
      		:uuid = "e5166dfd-81b7-3a4f-b993-ab68a010200d" ;
      		:version = "033" ;
      } // group ANC26-08

    group: ANC28 {

      // group attributes:
      		:description = "DTU Mean Sea Surface re-referenced to the WGS84 ellipsoid." ;
      		:fileName = "dtu13_20180705_001_01.nc" ;
      		:shortName = "ANC28" ;
      		:uuid = "56f47040-a72e-3109-99c2-bc1658e6dda4" ;
      		:version = "20180705" ;
      } // group ANC28

    group: ANC33 {

      // group attributes:
      		:description = "Water Mask File" ;
      		:fileName = "watermask_2000_20180301_001_global.h5" ;
      		:shortName = "ANC33" ;
      		:uuid = "1e7d3697-c576-308d-9197-21d827ac21db" ;
      		:version = "20180301" ;
      } // group ANC33

    group: ANC34 {

      // group attributes:
      		:description = "Urban Mask File" ;
      		:fileName = "SET_BY_PGE" ;
      		:shortName = "SET_BY_PGE" ;
      		:uuid = "SET_BY_PGE" ;
      		:version = "SET_BY_PGE" ;
      } // group ANC34

    group: ANC36-08 {

      // group attributes:
      		:description = "ISO 19139 XML file containing Series-level metadata information." ;
      		:fileName = "ATL08.003.series.xml" ;
      		:shortName = "ANC36-08" ;
      		:uuid = "a657d995-87c8-3a52-b4d4-d0de583b44ab" ;
      		:version = "003" ;
      } // group ANC36-08

    group: ANC38-08 {

      // group attributes:
      		:description = "ISO 19139 XML file containing DataSet-level metadata information." ;
      		:fileName = "ATL08.003.dataset.xml" ;
      		:shortName = "ANC38-08" ;
      		:uuid = "7ffd96d6-9c36-3ef7-80ab-606168059962" ;
      		:version = "003" ;
      } // group ANC38-08

    group: ATL03 {

      // group attributes:
      		:description = "ICESat-2 ATLAS L2A Global Geolocated Photon data products." ;
      		:fileName = "ATL03_20181014084920_02400109_003_01.h5" ;
      		:shortName = "ATL03" ;
      		:uuid = "498a71af-4c55-3685-bbe3-a704a1876765" ;
      		:version = "003" ;
      		:start_cycle = 1 ;
      		:end_cycle = 1 ;
      		:start_orbit = 441 ;
      		:end_orbit = 441 ;
      		:start_rgt = 240 ;
      		:end_rgt = 240 ;
      		:start_region = 9 ;
      		:end_region = 9 ;
      		:start_geoseg = 1151688 ;
      		:end_geoseg = 1280087 ;
      } // group ATL03

    group: ATL09 {

      // group attributes:
      		:description = "ICESat-2 ATLAS L3A atmosphere data products." ;
      		:fileName = "ATL09_20181014075514_02400101_003_01.h5" ;
      		:shortName = "ATL09" ;
      		:uuid = "ff8cd64b-f8d7-39e2-8b7f-f593d0477827" ;
      		:version = "003" ;
      		:start_cycle = 1 ;
      		:end_cycle = 1 ;
      		:start_orbit = 441 ;
      		:end_orbit = 441 ;
      		:start_rgt = 240 ;
      		:end_rgt = 240 ;
      		:start_region = 1 ;
      		:end_region = 14 ;
      		:start_geoseg = 12 ;
      		:end_geoseg = 2007117 ;
      } // group ATL09

    group: Control {

      // group attributes:
      		:description = "Text-based keyword=value file generated automatically within the ICESat-2 data system that specifies all of the conditions required for each individual run of the software." ;
      		:fileName = "CTL_atlas_l3a_ld_003713657.ctl" ;
      		:shortName = "CNTL" ;
      		:version = "1" ;
      } // group Control
    } // group Lineage

  group: ProcessStep {

    group: Browse {

      // group attributes:
      		:processDescription = "Browse processing is performed for each granule SIPS produces.  The browse utility reads data from the granule and produces browse images as defined in the respective product ATBD. The utility then embeds each browse image into the product within the /Browse group." ;
      		:identifier = "atlas_brw" ;
      		:softwareVersion = "Version 2.3" ;
      		:softwareDate = "Feb 14 2020" ;
      		:softwareTitle = "Creates ATLAS HDF5 browse files" ;
      		:runTimeParameters = "CTL_atlas_l3a_ld_003713657.ctl" ;
      		:stepDateTime = "2020-04-01T14:03:34.000000Z" ;
      } // group Browse

    group: Metadata {

      // group attributes:
      		:processDescription = "Metadata information is processed by the metadata utility for each granule produced by SIPS. During PGE processing, dynamic metadata are written to the product. Additional static information is provided with the metadata template. The metadata utility reads ISO Dataset and Series metadata files and updates the product with static information from within those files. The utility then merges the static and dynamic metadata to creates output ISO19139 Dataset and Series XML files. Finally the utility reads the ISO19139 Dataset and Series XML files into memory and stores the textual representations as attributes attached  to the /METADATA group." ;
      		:identifier = "atlas_meta" ;
      		:softwareVersion = "Version 4.3" ;
      		:softwareDate = "Feb  3 2020" ;
      		:softwareTitle = "Creates ATLAS XML metadata files" ;
      		:runTimeParameters = "CTL_atlas_l3a_ld_003713657.ctl" ;
      		:stepDateTime = "2020-04-01T14:03:36.000000Z" ;
      } // group Metadata

    group: PGE {

      // group attributes:
      		:ATBDDate = "01/17/2020" ;
      		:ATBDTitle = "Algorithm Theoretical Basis Document (ATBD) for Land - Vegetation Along-Track Products (ATL08)" ;
      		:ATBDVersion = "v.3" ;
      		:documentDate = "Feb 2020" ;
      		:documentation = "ATLAS Science Algorithm Software Design Description (SDD) - Volume 12 (atlas_l3a_ld)" ;
      		:processDescription = "Determines heights of ground and canopy surface. Where data permits, includes estimates of canopy height, relative canopy cover, canopy height distributions, surface roughness, surface slope/aspect and apparent reflectance." ;
      		:identifier = "atlas_l3a_ld" ;
      		:softwareVersion = "Version 3.3.1" ;
      		:softwareDate = "Mar 20 2020" ;
      		:softwareTitle = "ASAS L3A Land PGE" ;
      		:runTimeParameters = "CTL_atlas_l3a_ld_003713657.ctl" ;
      		:stepDateTime = "2020-04-01T14:03:26.000000Z" ;
      } // group PGE

    group: QA {

      // group attributes:
      		:processDescription = "QA processing is performed by an external utility on each granule produced by SIPS. The utility reads the granule, performs both generic and product-specific quality-assessment calculations, and writes a text-based quality assessment report. The name and creation data of this report are identified within the QADatasetIdentification metadata" ;
      		:identifier = "atl08_qa_util" ;
      		:softwareVersion = "Version 3.3" ;
      		:softwareDate = "Feb 14 2020" ;
      		:softwareTitle = "ATL08 QA Utility" ;
      		:runTimeParameters = "CTL_atlas_l3a_ld_003713657.ctl" ;
      		:stepDateTime = "2020-04-01T14:03:34.000000Z" ;
      } // group QA
    } // group ProcessStep

  group: ProductSpecificationDocument {

    // group attributes:
    		:ShortName = "ATL08_SDP" ;
    		:characterSet = "utf8" ;
    		:edition = "v4.3" ;
    		:language = "eng" ;
    		:publicationDate = "Feb 2020" ;
    		:title = "ICESat-2-SIPS-SPEC-4262 - ATLAS Science Algorithm Standard Data Product (SDP) Volume 7 (ATL08)." ;
    } // group ProductSpecificationDocument

  group: QADatasetIdentification {

    // group attributes:
    		:abstract = "An ASCII product that contains statistical information on data product results. These statistics enable data producers and users to assess the quality of the data in the data product granule" ;
    		:creationDate = "2020-04-01T14:03:34.000000Z" ;
    		:fileName = "ATL08_20181014084920_02400109_003_01.qa" ;
    } // group QADatasetIdentification

  group: SeriesIdentification {

    // group attributes:
    		:maintenanceAndUpdateFrequency = "asNeeded" ;
    		:maintenanceDate = "SET_BY_META" ;
    		:VersionID = "003" ;
    		:language = "eng" ;
    		:characterSet = "utf8" ;
    		:pointOfContact = "NSIDC DAAC > NASA National Snow and Ice Data Center Distributed Active Archive Center" ;
    		:longName = "ATLAS/ICESat-2 L3A Land and Vegetation Height" ;
    		:shortName = "ATL08" ;
    		:identifier_product_DOI = "doi:10.5067/ATLAS/ATL08.003" ;
    		:revisionDate = "2016-06-09" ;
    		:resourceProviderOrganizationName = "National Aeronautics and Space Administration (NASA)" ;
    		:abstract = "The ICESat-2 ATL08 standard data product contains along-track heights of ground and canopy surface at varying length scales. Where data permits, this includes estimates of canopy height, relative canopy cover, canopy height distributions, surface roughness, surface slope/aspect, and apparent reflectance." ;
    		:purpose = "The purpose of ATL08 is to provide along-track land/canopy heights and associated statistics." ;
    		:credit = "The software that generates the ATL08 product was designed and implemented within the ICESat-2 Science Investigator-led Processing System at the NASA Goddard Space Flight Center in Greenbelt, Maryland." ;
    		:status = "onGoing" ;
    		:format = "HDF" ;
    		:formatVersion = "5" ;
    		:topicCategory = "geoscientificInformation" ;
    		:mission = "ICESat-2 > Ice, Cloud, and land Elevation Satellite-2" ;
    } // group SeriesIdentification
  } // group METADATA

group: gt1r {

  // group attributes:
  		:Description = "Each group contains the segments for one Ground Track. As ICESat-2 orbits the earth, sequential transmit pulses illuminate six ground tracks on the surface of the earth.  The track width is approximately 14m.  Each ground track is numbered, according to the laser spot number that generates a given ground track.  Ground tracks are numbered from the left to the right in the direction of spacecraft travel as: 1L, 1R in the left-most pair of beams; 2L, 2R for the center pair of beams; and 3L, 3R for the right-most pair of beams." ;
  		:atlas_pce = "pce3" ;
  		:atlas_beam_type = "strong" ;
  		:groundtrack_id = "gt1r" ;
  		:atmosphere_profile = "profile_1" ;
  		:atlas_spot_number = "5" ;
  		:sc_orientation = "Forward" ;

  group: signal_photons {
    dimensions:
    	delta_time = UNLIMITED ; // (1185 currently)
    variables:
    	byte classed_pc_flag(delta_time) ;
    		classed_pc_flag:coordinates = "delta_time" ;
    		classed_pc_flag:description = "Land Vegetation ATBD classification flag for each photon as either noise, ground, canopy, and top of canopy. 0 = noise,  1 = ground, 2 = canopy, or 3 = top of canopy." ;
    		classed_pc_flag:flag_meanings = "noise ground canopy top_of_canopy" ;
    		classed_pc_flag:flag_values = 0b, 1b, 2b, 3b ;
    		classed_pc_flag:long_name = "photon land atbd classification" ;
    		classed_pc_flag:source = "Land ATBD section 4.10" ;
    		classed_pc_flag:units = "1" ;
    	int classed_pc_indx(delta_time) ;
    		classed_pc_indx:contentType = "referenceInformation" ;
    		classed_pc_indx:coordinates = "delta_time" ;
    		classed_pc_indx:description = "Index  (1-based) of the ATL08 classified signal photon from the start of the ATL03 geolocation segment specified on the ATL08 product at the photon rate in the corresponding parameter, ph_segment_id. This index traces back to specific photon within a 20m segment_id on ATL03.  The unique identifier for tracing each ATL08 signal photon to the corresponding photon record on ATL03 is the segment_id, orbit, cycle, and classed_pc_indx. Orbit and cycle intervals for the granule are found in the /ancillary_data. The timestamp of each orbit transition is found in the /orbit_info group." ;
    		classed_pc_indx:long_name = "indicies of classed photons" ;
    		classed_pc_indx:source = "Retained from prior a_alt_science_ph packet" ;
    		classed_pc_indx:units = "1" ;
    	byte d_flag(delta_time) ;
    		d_flag:coordinates = "delta_time" ;
    		d_flag:description = "Flag indicating the labeling of DRAGANN noise filtering for a given photon." ;
    		d_flag:flag_meanings = "noise signal" ;
    		d_flag:flag_values = 0b, 1b ;
    		d_flag:long_name = "dragann flag" ;
    		d_flag:source = "Land ATBD section 2.3.5" ;
    		d_flag:units = "1" ;
    	double delta_time(delta_time) ;
    		delta_time:description = "Number of GPS seconds since the ATLAS SDP epoch. The ATLAS Standard Data Products (SDP) epoch offset is defined within /ancillary_data/atlas_sdp_gps_epoch as the number of GPS seconds between the GPS epoch (1980-01-06T00:00:00.000000Z UTC) and the ATLAS SDP epoch. By adding the offset contained within atlas_sdp_gps_epoch to delta time parameters, the time in gps_seconds relative to the GPS epoch can be computed." ;
    		delta_time:long_name = "delta time" ;
    		delta_time:source = "ATL03" ;
    		delta_time:standard_name = "time" ;
    		delta_time:units = "seconds since 2018-01-01" ;
    	int ph_segment_id(delta_time) ;
    		ph_segment_id:contentType = "referenceInformation" ;
    		ph_segment_id:coordinates = "delta_time" ;
    		ph_segment_id:description = "Segment ID of photons tracing back to specific 20m segment_id on ATL03.  The unique identifier for tracing each ATL08 signal photon to the photon on ATL03 is the segment_id, orbit, and classed_pc_indx. The unique identifier for tracing each ATL08 signal photon to the corresponding photon record on ATL03 is the segment_id, orbit, cycle, and classed_pc_indx. Orbit and cycle intervals for the granule are found in the /ancillary_data. The timestamp of each orbit transition is found in the /orbit_info group." ;
    		ph_segment_id:long_name = "segment id of photon" ;
    		ph_segment_id:source = "Retained from prior a_alt_science_ph packet" ;
    		ph_segment_id:units = "1" ;

    // group attributes:
    		:Description = "Contains parameters related to individual photons." ;
    		:data_rate = "Data are stored at the signal-photon classification rate." ;
    } // group signal_photons

  group: land_segments {
    dimensions:
    	delta_time = UNLIMITED ; // (5 currently)
    variables:
    	float asr(delta_time) ;
    		asr:_FillValue = 3.402823e+38f ;
    		asr:coordinates = "delta_time latitude longitude" ;
    		asr:description = "Apparent surface reflectance" ;
    		asr:long_name = "apparent surface reflectance" ;
    		asr:source = "ATL09" ;
    		asr:units = "1" ;
    	float atlas_pa(delta_time) ;
    		atlas_pa:_FillValue = 3.402823e+38f ;
    		atlas_pa:contentType = "referenceInformation" ;
    		atlas_pa:coordinates = "delta_time latitude longitude" ;
    		atlas_pa:description = "Off nadir pointing angle (in radians) of the satellite to increase spatial sampling in the non-polar regions. ATLAS_PA =90degs-beam_coelev." ;
    		atlas_pa:long_name = "atlas pointing angle" ;
    		atlas_pa:source = "ATL03" ;
    		atlas_pa:units = "radians" ;
    	float beam_azimuth(delta_time) ;
    		beam_azimuth:_FillValue = 3.402823e+38f ;
    		beam_azimuth:contentType = "referenceInformation" ;
    		beam_azimuth:coordinates = "delta_time latitude longitude" ;
    		beam_azimuth:description = "Azimuth(in radians) of the unit pointing vector for the reference photon in the local ENU frame in radians.  The angle is measured from north and positive towards East." ;
    		beam_azimuth:long_name = "beam azimuth" ;
    		beam_azimuth:source = "ATL03" ;
    		beam_azimuth:units = "radians" ;
    	float beam_coelev(delta_time) ;
    		beam_coelev:_FillValue = 3.402823e+38f ;
    		beam_coelev:contentType = "referenceInformation" ;
    		beam_coelev:coordinates = "delta_time latitude longitude" ;
    		beam_coelev:description = "Co-elevation (CE) is direction from vertical of the laser beam as seen by an observer located at the laser ground spot." ;
    		beam_coelev:long_name = "beam co-elevation" ;
    		beam_coelev:source = "ATL03" ;
    		beam_coelev:units = "radians" ;
    	byte brightness_flag(delta_time) ;
    		brightness_flag:_FillValue = 127b ;
    		brightness_flag:coordinates = "delta_time latitude longitude" ;
    		brightness_flag:description = "Flag indicating that the ground surface is bright (e.g. snow-covered or other bright surfaces)" ;
    		brightness_flag:flag_meanings = "not_bright_surface bright_surface" ;
    		brightness_flag:flag_values = 0b, 1b ;
    		brightness_flag:long_name = "brightness flag" ;
    		brightness_flag:source = "Land ATBD section 2.4.21" ;
    		brightness_flag:units = "1" ;
    	byte cloud_flag_atm(delta_time) ;
    		cloud_flag_atm:_FillValue = 127b ;
    		cloud_flag_atm:coordinates = "delta_time latitude longitude" ;
    		cloud_flag_atm:description = "Cloud confidence flag from ATL09 that indicates the number of cloud or aerosol layers identified in each 25Hz atmospheric profile. If the flag is greater than 0, aerosols or clouds could be present. Valid range is 0 - 10." ;
    		cloud_flag_atm:long_name = "cloud flag atm" ;
    		cloud_flag_atm:source = "ATL09" ;
    		cloud_flag_atm:units = "1" ;
    		cloud_flag_atm:valid_max = 10b ;
    		cloud_flag_atm:valid_min = 0b ;
    	byte cloud_fold_flag(delta_time) ;
    		cloud_fold_flag:coordinates = "delta_time latitude longitude" ;
    		cloud_fold_flag:description = "Flag that indicates this profile likely contains cloud signal folded down from above 15 km to the last 2-3 km of the profile. See ATL09 ATBD Table 3.9 for detailed flag value meanings." ;
    		cloud_fold_flag:flag_meanings = "no_folding goes5_indicates profile_indicates both_indicate" ;
    		cloud_fold_flag:flag_values = 0b, 1b, 2b, 3b ;
    		cloud_fold_flag:long_name = "cloud folding flag" ;
    		cloud_fold_flag:source = "ATL09" ;
    		cloud_fold_flag:valid_max = 3b ;
    		cloud_fold_flag:valid_min = 0b ;
    		cloud_fold_flag:_FillValue = 127b ;
    		cloud_fold_flag:contentType = "modelResult" ;
    	double delta_time(delta_time) ;
    		delta_time:coordinates = "latitude longitude" ;
    		delta_time:description = "Mean time for the segment in number of GPS seconds since the ATLAS SDP epoch. The ATLAS Standard Data Products (SDP) epoch offset is defined within /ancillary_data/atlas_sdp_gps_epoch as the number of GPS seconds between the GPS epoch (1980-01-06T00:00:00.000000Z UTC) and the ATLAS SDP epoch. By adding the offset contained within atlas_sdp_gps_epoch to delta time parameters, the time in gps_seconds relative to the GPS epoch can be computed." ;
    		delta_time:long_name = "mean_pass_time" ;
    		delta_time:source = "Land ATBD section 2.4" ;
    		delta_time:standard_name = "time" ;
    		delta_time:units = "seconds since 2018-01-01" ;
    	double delta_time_beg(delta_time) ;
    		delta_time_beg:contentType = "referenceInformation" ;
    		delta_time_beg:coordinates = "delta_time latitude longitude" ;
    		delta_time_beg:description = "Time of the first photon contained within the data segment, in seconds since the ATLAS SDP GPS Epoch. The ATLAS Standard Data Products (SDP) epoch offset is defined within /ancillary_data/atlas_sdp_gps_epoch as the number of GPS seconds between the GPS epoch (1980-01-06T00:00:00.000000Z UTC) and the ATLAS SDP epoch. By adding the offset contained within atlas_sdp_gps_epoch to delta time parameters, the time in gps_seconds relative to the GPS epoch can be computed." ;
    		delta_time_beg:long_name = "delta time begin" ;
    		delta_time_beg:source = "Derived (gps_seconds-gps_sec_offset)" ;
    		delta_time_beg:units = "seconds since 2018-01-01" ;
    	double delta_time_end(delta_time) ;
    		delta_time_end:contentType = "referenceInformation" ;
    		delta_time_end:coordinates = "delta_time latitude longitude" ;
    		delta_time_end:description = "Time of the last photon contained within the data segment, in seconds since the ATLAS SDP epoch. The ATLAS Standard Data Products (SDP) epoch offset is defined within /ancillary_data/atlas_sdp_gps_epoch as the number of GPS seconds between the GPS epoch (1980-01-06T00:00:00.000000Z UTC) and the ATLAS SDP epoch. By adding the offset contained within atlas_sdp_gps_epoch to delta time parameters, the time in gps_seconds relative to the GPS epoch can be computed." ;
    		delta_time_end:long_name = "delta time end" ;
    		delta_time_end:source = "Derived (gps_seconds-gps_sec_offset)" ;
    		delta_time_end:units = "seconds since 2018-01-01" ;
    	byte dem_flag(delta_time) ;
    		dem_flag:_FillValue = 127b ;
    		dem_flag:contentType = "referenceInformation" ;
    		dem_flag:coordinates = "delta_time latitude longitude" ;
    		dem_flag:description = "Indicates source of the DEM height. Values: 0=None, 1=Arctic, 2=GMTED, 3=MSS, 4=Antarctic." ;
    		dem_flag:flag_meanings = "none arctic gmted mss antarctic" ;
    		dem_flag:flag_values = 0b, 1b, 2b, 3b, 4b ;
    		dem_flag:long_name = "dem source flag" ;
    		dem_flag:source = "Atmosphere ATBD" ;
    		dem_flag:units = "1" ;
    		dem_flag:valid_max = 4b ;
    		dem_flag:valid_min = 0b ;
    	float dem_h(delta_time) ;
    		dem_h:_FillValue = 3.402823e+38f ;
    		dem_h:contentType = "referenceInformation" ;
    		dem_h:coordinates = "delta_time latitude longitude" ;
    		dem_h:description = "Best available DEM (in priority of Arctic/Antarctic/GMTED/MSS) value at the geolocation point.  Height is in meters above the WGS84 Ellipsoid." ;
    		dem_h:long_name = "dem height" ;
    		dem_h:source = "GIMP, GMTED,MSS" ;
    		dem_h:units = "meters" ;
    	byte dem_removal_flag(delta_time) ;
    		dem_removal_flag:coordinates = "delta_time latitude longitude" ;
    		dem_removal_flag:description = "Flag indicating more than dem_removal_percent_limit (default 20.0) removed from land segment due to failing DEM-QA tests" ;
    		dem_removal_flag:flag_meanings = "below_threshold above_threshold" ;
    		dem_removal_flag:flag_values = 0b, 1b ;
    		dem_removal_flag:long_name = "dem removal flag" ;
    		dem_removal_flag:source = "ATBD section 2.4.11" ;
    		dem_removal_flag:units = "1" ;
    	float h_dif_ref(delta_time) ;
    		h_dif_ref:_FillValue = 3.402823e+38f ;
    		h_dif_ref:coordinates = "delta_time latitude longitude" ;
    		h_dif_ref:description = "Difference between h_te_median and ref_DEM" ;
    		h_dif_ref:long_name = "h dif from reference" ;
    		h_dif_ref:source = "Land ATBD section 2.4" ;
    		h_dif_ref:units = "meters" ;
    	float last_seg_extend(delta_time) ;
    		last_seg_extend:coordinates = "delta_time latitude longitude" ;
    		last_seg_extend:description = "The distance (km) that the last ATL08 processing segment in a file is either extended or overlapped with the previous ATL08 processing segment." ;
    		last_seg_extend:long_name = "last segment extended" ;
    		last_seg_extend:source = "Land ATBD 13March2019, Section 2.4.20" ;
    		last_seg_extend:standard_name = "last_seg_extend" ;
    		last_seg_extend:units = "kilometers" ;
    	float latitude(delta_time) ;
    		latitude:coordinates = "delta_time longitude" ;
    		latitude:description = "Latitude of the center-most signal photon within each segment." ;
    		latitude:long_name = "latitude" ;
    		latitude:source = "Land ATBD section 2.4" ;
    		latitude:standard_name = "latitude" ;
    		latitude:units = "degrees" ;
    		latitude:valid_max = 90.f ;
    		latitude:valid_min = -90.f ;
    	byte layer_flag(delta_time) ;
    		layer_flag:contentType = "modelResult" ;
    		layer_flag:coordinates = "delta_time latitude longitude" ;
    		layer_flag:description = "This flag is a combination of multiple flags (cloud_flag_atm, cloud_flag_asr, and bsnow_con) and takes daytime/nighttime into consideration. A value of 1 means clouds or blowing snow are likely present. A value of 0 indicates the likely absence of clouds or blowing snow." ;
    		layer_flag:flag_meanings = "likely_clear likely_cloudy" ;
    		layer_flag:flag_values = 0b, 1b ;
    		layer_flag:long_name = "consolidated cloud flag" ;
    		layer_flag:source = "ATL09" ;
    	float longitude(delta_time) ;
    		longitude:coordinates = "delta_time latitude" ;
    		longitude:description = "Longitude of the center-most signal photon within each segment." ;
    		longitude:long_name = "longitude" ;
    		longitude:source = "Land ATBD section 2.4" ;
    		longitude:standard_name = "longitude" ;
    		longitude:units = "degrees" ;
    		longitude:valid_max = 180.f ;
    		longitude:valid_min = -180.f ;
    	byte msw_flag(delta_time) ;
    		msw_flag:_FillValue = 127b ;
    		msw_flag:coordinates = "delta_time latitude longitude" ;
    		msw_flag:description = "Multiple Scattering warning flag. The multiple scattering warning flag (ATL09 parameter msw_flag) has values from -1 to 5 where zero means no multiple scattering and 5 the greatest. If no layers were detected, then msw_flag = 0. If blowing snow is detected and its estimated optical depth is greater than or equal to 0.5, then msw_flag = 5. If the blowing snow optical depth is less than 0.5, then msw_flag = 4. If no blowing snow is detected but there are cloud or aerosol layers detected, the msw_flag assumes values of 1 to 3 based on the height of the bottom of the lowest layer: < 1 km, msw_flag = 3; 1-3 km, msw_flag = 2; > 3km, msw_flag = 1. A value of -1 indicates that the signal to noise of the data was too low to reliably ascertain the presence of cloud or blowing snow. We expect values of -1 to occur only during daylight." ;
    		msw_flag:flag_meanings = "cannot_determine no_layers layer_gt_3km layer_between_1_and_3_km layer_lt_1km blow_snow_od_lt_0.5 blow_snow_od_gt_0.5" ;
    		msw_flag:flag_values = -1b, 0b, 1b, 2b, 3b, 4b, 5b ;
    		msw_flag:long_name = "multiple scattering warning flag" ;
    		msw_flag:source = "ATL09" ;
    		msw_flag:units = "1" ;
    	int n_seg_ph(delta_time) ;
    		n_seg_ph:coordinates = "delta_time latitude longitude" ;
    		n_seg_ph:description = "Number of photons within each land segment." ;
    		n_seg_ph:long_name = "number of photons" ;
    		n_seg_ph:source = "Derived" ;
    		n_seg_ph:units = "1" ;
    	int night_flag(delta_time) ;
    		night_flag:_FillValue = 2147483647 ;
    		night_flag:coordinates = "delta_time latitude longitude" ;
    		night_flag:description = "Flag indicating the data were acquired in night conditions: 0=day, 1=night.  Flag is derived from solar elevation at the geolocated segment.  IF solar elevation is above threshold it is day, if not then it is night.  Threshold is set in atlas_l3a_const_mod." ;
    		night_flag:flag_meanings = "day night" ;
    		night_flag:flag_values = 0, 1 ;
    		night_flag:long_name = "night flag" ;
    		night_flag:source = "Land ATBD section 2.4.8" ;
    		night_flag:units = "1" ;
    	int64 ph_ndx_beg(delta_time) ;
    		ph_ndx_beg:coordinates = "delta_time latitude longitude" ;
    		ph_ndx_beg:description = "Index (1-based) within the photon-rate data (/land_segments/photons) of the first photon within this each land segment." ;
    		ph_ndx_beg:long_name = "photon index begin" ;
    		ph_ndx_beg:source = "Derived" ;
    		ph_ndx_beg:units = "1" ;
    	byte ph_removal_flag(delta_time) ;
    		ph_removal_flag:coordinates = "delta_time latitude longitude" ;
    		ph_removal_flag:description = "Flag indicating more than ph_removal_percent_limit (default 50.0) removed from land segment due to failing QA tests" ;
    		ph_removal_flag:flag_meanings = "below_threshold above_threshold" ;
    		ph_removal_flag:flag_values = 0b, 1b ;
    		ph_removal_flag:long_name = "ph removal flag" ;
    		ph_removal_flag:source = "ATBD section 4.13" ;
    		ph_removal_flag:units = "1" ;
    	byte psf_flag(delta_time) ;
    		psf_flag:contentType = "referenceInformation" ;
    		psf_flag:coordinates = "delta_time latitude longitude" ;
    		psf_flag:description = "Flag is set to 1 if the point spread function (computed as sigma_atlas_land) has exceeded the threshold (1 m)" ;
    		psf_flag:flag_meanings = "below_threshold above_threshold" ;
    		psf_flag:flag_values = 0b, 1b ;
    		psf_flag:long_name = "point spread function flag" ;
    		psf_flag:source = "Land/Veg ATBD" ;
    		psf_flag:units = "1" ;
    		psf_flag:valid_max = 1b ;
    		psf_flag:valid_min = 0b ;
    	short rgt(delta_time) ;
    		rgt:contentType = "referenceInformation" ;
    		rgt:coordinates = "delta_time latitude longitude" ;
    		rgt:description = "The reference ground track (RGT) is the track on the earth at which a specified unit vector within the observatory is pointed. Under nominal operating conditions, there will be no data collected along the RGT, as the RGT is spanned by GT3 and GT4.  During slews or off-pointing, it is possible that ground tracks may intersect the RGT. The ICESat-2 mission has 1387 RGTs." ;
    		rgt:long_name = "reference ground track" ;
    		rgt:source = "Operations" ;
    		rgt:units = "1" ;
    		rgt:valid_max = 1387s ;
    		rgt:valid_min = 1s ;
    	int segment_id_beg(delta_time) ;
    		segment_id_beg:contentType = "referenceInformation" ;
    		segment_id_beg:coordinates = "delta_time latitude longitude" ;
    		segment_id_beg:description = "Geolocation segment number of the first photon in the land segment." ;
    		segment_id_beg:long_name = "begin geolocation segment bin" ;
    		segment_id_beg:source = "ATL03" ;
    		segment_id_beg:units = "1" ;
    	int segment_id_end(delta_time) ;
    		segment_id_end:contentType = "referenceInformation" ;
    		segment_id_end:coordinates = "delta_time latitude longitude" ;
    		segment_id_end:description = "Geolocation segment number of the last photon in the land segment." ;
    		segment_id_end:long_name = "end geolocation segment bin" ;
    		segment_id_end:source = "ATL03" ;
    		segment_id_end:units = "1" ;
    	int segment_landcover(delta_time) ;
    		segment_landcover:_FillValue = 255 ;
    		segment_landcover:coordinates = "delta_time latitude longitude" ;
    		segment_landcover:description = "IGBP Land Cover Surface type classification as reference from MODIS Land Cover(ANC18) at the 0.5 arcsecond resolution." ;
    		segment_landcover:flag_meanings = "Water Evergreen_Needleleaf_Forest Evergreen_Broadleaf_Forest Deciduous_Needleleaf_Forest Deciduous_Broadleaf_Forest Mixed_Forest Closed_Shrublands Open_Shrubland Woody_Savanna Savanna Grassland Wetland Croplands Urban Crop_Mosaic Permanent_Snow Barren" ;
    		segment_landcover:flag_values = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16 ;
    		segment_landcover:long_name = "segment landcover" ;
    		segment_landcover:source = "ATBD section 2.4.14" ;
    		segment_landcover:units = "1" ;
    		segment_landcover:valid_max = 16 ;
    		segment_landcover:valid_min = 0 ;
    	byte segment_snowcover(delta_time) ;
    		segment_snowcover:_FillValue = 127b ;
    		segment_snowcover:coordinates = "delta_time latitude longitude" ;
    		segment_snowcover:description = "Daily snow/ice cover from ATL09 at the 25 Hz rate(275m) indicating likely presence of snow and ice within each segment. 0=ice free water; 1=snow free land;  2=snow; 3=ice." ;
    		segment_snowcover:flag_meanings = "ice_free_water snow_free_land snow ice" ;
    		segment_snowcover:flag_values = 0b, 1b, 2b, 3b ;
    		segment_snowcover:long_name = "segment snowcover" ;
    		segment_snowcover:source = "ATBD section 4.2.16" ;
    		segment_snowcover:units = "1" ;
    		segment_snowcover:valid_max = 3b ;
    		segment_snowcover:valid_min = 0b ;
    	int segment_watermask(delta_time) ;
    		segment_watermask:_FillValue = 255 ;
    		segment_watermask:coordinates = "delta_time latitude longitude" ;
    		segment_watermask:description = "Water mask(i.e. flag) indicating inland water as referenced from the Global Raster Water Mask(ANC33) at 250 m spatial resolution." ;
    		segment_watermask:flag_meanings = "no_water water" ;
    		segment_watermask:flag_values = 0, 1 ;
    		segment_watermask:long_name = "segment watermask" ;
    		segment_watermask:source = "ATBD section 2.4.15" ;
    		segment_watermask:units = "1" ;
    		segment_watermask:valid_max = 1 ;
    		segment_watermask:valid_min = 0 ;
    	float sigma_across(delta_time) ;
    		sigma_across:_FillValue = 3.402823e+38f ;
    		sigma_across:contentType = "referenceInformation" ;
    		sigma_across:coordinates = "delta_time latitude longitude" ;
    		sigma_across:description = "Total cross-track uncertainty due to PPD and POD knowledge.  Read from ATL03 product gtx/geolocation/sigma_across. Sigma_atlas_y is reported on ATL08 as the uncertainty of the center-most reference photon of the 100m ATL08 segment." ;
    		sigma_across:long_name = "sigma atlas y" ;
    		sigma_across:source = "ATL03" ;
    		sigma_across:units = "1" ;
    	float sigma_along(delta_time) ;
    		sigma_along:_FillValue = 3.402823e+38f ;
    		sigma_along:contentType = "referenceInformation" ;
    		sigma_along:coordinates = "delta_time latitude longitude" ;
    		sigma_along:description = "Total along-track uncertainty due to PPD and POD knowledge.  Read from ATL03 product gtx/geolocation/sigma_along. Sigma_atlas_x is reported on ATL08 as the uncertainty of the center-most reference photon of the 100m ATL08 segment." ;
    		sigma_along:long_name = "sigma atlas x" ;
    		sigma_along:source = "ATL03" ;
    		sigma_along:units = "1" ;
    	float sigma_atlas_land(delta_time) ;
    		sigma_atlas_land:_FillValue = 3.402823e+38f ;
    		sigma_atlas_land:contentType = "referenceInformation" ;
    		sigma_atlas_land:coordinates = "delta_time latitude longitude" ;
    		sigma_atlas_land:description = "Total vertical geolocation error due to ranging and local surface slope.  The parameter is computed for ATL08 as described in equation 1.2." ;
    		sigma_atlas_land:long_name = "sigma atlas land" ;
    		sigma_atlas_land:source = "Land ATBD section 2.5.13" ;
    		sigma_atlas_land:units = "1" ;
    	float sigma_h(delta_time) ;
    		sigma_h:_FillValue = 3.402823e+38f ;
    		sigma_h:contentType = "referenceInformation" ;
    		sigma_h:coordinates = "delta_time latitude longitude" ;
    		sigma_h:description = "Estimated uncertainty for the reference photon bounce point ellipsoid height: 1- sigma (m) provided at the geolocation segment rate on ATL03.  Sigma_h is reported on ATL08 as the uncertainty of the center-most reference photon of the 100m ATL08 segment." ;
    		sigma_h:long_name = "height uncertainty" ;
    		sigma_h:source = "ATL03" ;
    		sigma_h:units = "1" ;
    	float sigma_topo(delta_time) ;
    		sigma_topo:_FillValue = 3.402823e+38f ;
    		sigma_topo:contentType = "referenceInformation" ;
    		sigma_topo:coordinates = "delta_time latitude longitude" ;
    		sigma_topo:description = "Total uncertainty that include sigma_h plus geolocation uncertainty due to local slope (equation 1.3).  The local slope is multiplied by the geolocation uncertainty factor. This will be used to determine the total vertical geolocation error due to ranging and local slope." ;
    		sigma_topo:long_name = "sigma atlas topo" ;
    		sigma_topo:source = "Land ATBD section 2.5.12" ;
    		sigma_topo:units = "1" ;
    	float snr(delta_time) ;
    		snr:_FillValue = 3.402823e+38f ;
    		snr:coordinates = "delta_time latitude longitude" ;
    		snr:description = "The signal to noise ratio of geolocated photons as determined by the ratio of the superset of ATL03 signal and DRAGANN found signal photons used for processing the ATL08 segments to the background photons (i.e. noise) within the same ATL08 segments." ;
    		snr:long_name = "signal to noise ratio" ;
    		snr:source = "ATBD section 2.5.14" ;
    		snr:units = "1" ;
    	float solar_azimuth(delta_time) ;
    		solar_azimuth:contentType = "referenceInformation" ;
    		solar_azimuth:coordinates = "delta_time latitude longitude" ;
    		solar_azimuth:description = "The direction, eastwards from north, of the sun vector as seen by an observer at the laser ground spot." ;
    		solar_azimuth:long_name = "solar azimuth" ;
    		solar_azimuth:source = "ATL03g ATBD" ;
    		solar_azimuth:units = "degrees_east" ;
    	float solar_elevation(delta_time) ;
    		solar_elevation:contentType = "referenceInformation" ;
    		solar_elevation:coordinates = "delta_time latitude longitude" ;
    		solar_elevation:description = "Solar Angle above or below the plane tangent to the ellipsoid surface at the laser spot. Positive values mean the sun is above the horizon, while  negative values mean it is below the horizon. The effect of atmospheric refraction is not included. This is a low precision value, with approximately TBD degree accuracy." ;
    		solar_elevation:long_name = "solar elevation" ;
    		solar_elevation:source = "ATL03g ATBD" ;
    		solar_elevation:units = "degrees" ;
    	byte surf_type(delta_time, ds_surf_type) ;
    		surf_type:contentType = "referenceInformation" ;
    		surf_type:coordinates = "delta_time latitude longitude" ;
    		surf_type:description = "Flags describing which surface types this interval is associated with. 0=not type, 1=is type. Order of array is land, ocean, sea ice, land ice, inland water." ;
    		surf_type:flag_meanings = "not_type is_type" ;
    		surf_type:flag_values = 0b, 1b ;
    		surf_type:long_name = "surface type" ;
    		surf_type:source = "ATL03 ATBD, Section 4" ;
    		surf_type:units = "1" ;
    		surf_type:valid_max = 1b ;
    		surf_type:valid_min = 0b ;
    	int terrain_flg(delta_time) ;
    		terrain_flg:_FillValue = 2147483647 ;
    		terrain_flg:coordinates = "delta_time latitude longitude" ;
    		terrain_flg:description = "Terrain flag quality check to indicate a deviation above a threshold from the reference DEM height reported on the product." ;
    		terrain_flg:flag_meanings = "below_threshold above_threshold" ;
    		terrain_flg:flag_values = 0, 1 ;
    		terrain_flg:long_name = "terrain flag" ;
    		terrain_flg:source = "Land ATBD section 2.4.8" ;
    		terrain_flg:units = "1" ;
    	int urban_flag(delta_time) ;
    		urban_flag:_FillValue = 2147483647 ;
    		urban_flag:coordinates = "delta_time latitude longitude" ;
    		urban_flag:description = "The urban flag indicates that a segment is likely located over an urban area." ;
    		urban_flag:flag_meanings = "not_urban urban" ;
    		urban_flag:flag_values = 0, 1 ;
    		urban_flag:long_name = "segment urban flag" ;
    		urban_flag:source = "Land ATBD section 2.4.17" ;
    		urban_flag:units = "1" ;

    // group attributes:
    		:Description = "Contains data categorized as land at 100 meter intervals." ;
    		:data_rate = "Data are stored as aggregates of 100 meters." ;

    group: canopy {
      variables:
      	int canopy_flag(delta_time) ;
      		canopy_flag:_FillValue = 2147483647 ;
      		canopy_flag:coordinates = "../delta_time ../latitude ../longitude" ;
      		canopy_flag:description = "Flag indicating that canopy was detected using the Landsat Tree Cover Continuous Fields data product. If percent of canopy cover along the L-km segment is greater than 5%, then canopy is assumed to be present; else, no canopy is assumed present." ;
      		canopy_flag:flag_meanings = "no_canopy_present canopy_present" ;
      		canopy_flag:flag_values = 0, 1 ;
      		canopy_flag:long_name = "canopy flag" ;
      		canopy_flag:source = "Land ATBD section 2.2.22" ;
      		canopy_flag:units = "1" ;
      	float canopy_h_metrics(delta_time, ds_metrics) ;
      		canopy_h_metrics:_FillValue = 3.402823e+38f ;
      		canopy_h_metrics:coordinates = "../delta_time ../latitude ../longitude" ;
      		canopy_h_metrics:description = "Height metrics based on the cumulative distribution of relative canopy heights above the interpolated ground surface.  The height metrics are calculated at the following percentiles: 25,50,60,70,75,80,85,90,95%." ;
      		canopy_h_metrics:long_name = "canopy height metrics" ;
      		canopy_h_metrics:source = "Land ATBD section 2.2.3" ;
      		canopy_h_metrics:units = "meters" ;
      	float canopy_h_metrics_abs(delta_time, ds_metrics) ;
      		canopy_h_metrics_abs:_FillValue = 3.402823e+38f ;
      		canopy_h_metrics_abs:coordinates = "../delta_time ../latitude ../longitude" ;
      		canopy_h_metrics_abs:description = "Height metrics based on the cumulative distribution of absolute canopy heights above the WGS84 Ellipsoid.  The height metrics are calculated at the following percentiles: 25,50,60,70,75,80,85,90,95%." ;
      		canopy_h_metrics_abs:long_name = "canopy absolute height metrics" ;
      		canopy_h_metrics_abs:source = "Land ATBD section 2.2.3" ;
      		canopy_h_metrics_abs:units = "meters" ;
      	float canopy_openness(delta_time) ;
      		canopy_openness:_FillValue = 3.402823e+38f ;
      		canopy_openness:coordinates = "../delta_time ../latitude ../longitude" ;
      		canopy_openness:description = "Standard Deviation of all photons classified as canopy photons within the segment to provide inference of canopy openness." ;
      		canopy_openness:long_name = "canopy openness" ;
      		canopy_openness:source = "Land ATBD section 4.12" ;
      		canopy_openness:units = "1" ;
      	byte canopy_rh_conf(delta_time) ;
      		canopy_rh_conf:contentType = "modelResult" ;
      		canopy_rh_conf:coordinates = "../delta_time ../latitude ../longitude" ;
      		canopy_rh_conf:description = "Canopy relative height confidence flag based on percentage of ground and canopy photons within a segment: 0 (<5% canopy), 1 (>5% canopy, <5% ground), 2 (>5% canopy, >5% ground)." ;
      		canopy_rh_conf:flag_meanings = "<5%_canopy >=5%_canopy_<5%_ground >=5%_canopy_>=5%_ground" ;
      		canopy_rh_conf:flag_values = 0b, 1b, 2b ;
      		canopy_rh_conf:long_name = "canopy relative height confidence" ;
      		canopy_rh_conf:source = "Land/Veg ATBD 13March2019, Section 2.2.21" ;
      		canopy_rh_conf:units = "1" ;
      		canopy_rh_conf:valid_max = 2b ;
      		canopy_rh_conf:valid_min = 0b ;
      	float centroid_height(delta_time) ;
      		centroid_height:_FillValue = 3.402823e+38f ;
      		centroid_height:coordinates = "../delta_time ../latitude ../longitude" ;
      		centroid_height:description = "Optical centroid of all photons classified as either canopy or ground points within the segment.  The heights used in this calculation are absolute heights above the reference ellipsoid. This parameter is equivalent to the centroid height produced ICESat GLA14." ;
      		centroid_height:long_name = "centroid height" ;
      		centroid_height:source = "Land ATBD section 2.2.22" ;
      		centroid_height:units = "meters" ;
      	float h_canopy(delta_time) ;
      		h_canopy:_FillValue = 3.402823e+38f ;
      		h_canopy:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_canopy:description = "98% height of all the individual canopy relative heights for the segment above the estimated terrain surface. Relative canopy heights have been computed by differencing the canopy photon height from the estimated terrain surface." ;
      		h_canopy:long_name = "height canopy" ;
      		h_canopy:source = "Land ATBD section 4.12" ;
      		h_canopy:units = "meters" ;
      	float h_canopy_abs(delta_time) ;
      		h_canopy_abs:_FillValue = 3.402823e+38f ;
      		h_canopy_abs:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_canopy_abs:description = "The 98% height of all the absolute individual canopy heights referenced above the WGS84 ellipsoid." ;
      		h_canopy_abs:long_name = "absolute segment canopy height" ;
      		h_canopy_abs:source = "Land ATBD section 2.2.2" ;
      		h_canopy_abs:units = "meters" ;
      	float h_canopy_quad(delta_time) ;
      		h_canopy_quad:_FillValue = 3.402823e+38f ;
      		h_canopy_quad:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_canopy_quad:description = "The quadratic mean height of individual classified relative canopy photon heights above the estimated terrain surface." ;
      		h_canopy_quad:long_name = "canopy quadratic mean" ;
      		h_canopy_quad:source = "Land ATBD section 4.12" ;
      		h_canopy_quad:units = "meters" ;
      	float h_canopy_uncertainty(delta_time) ;
      		h_canopy_uncertainty:_FillValue = 3.402823e+38f ;
      		h_canopy_uncertainty:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_canopy_uncertainty:description = "Uncertainty of the relative canopy heights for the segment. Incorporates all systematic uncertainties as well as uncertainty from errors of identified photons. See section 1 and equations 1.4 and 1.5 in the Land ATBD" ;
      		h_canopy_uncertainty:long_name = "segment canopy height uncertainty" ;
      		h_canopy_uncertainty:source = "Land ATBD section 1.5" ;
      		h_canopy_uncertainty:units = "meters" ;
      	float h_dif_canopy(delta_time) ;
      		h_dif_canopy:_FillValue = 3.402823e+38f ;
      		h_dif_canopy:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_dif_canopy:description = "Difference between h_canopy and h_median_canopy" ;
      		h_dif_canopy:long_name = "canopy diff to median height" ;
      		h_dif_canopy:source = "Land ATBD section 4.12" ;
      		h_dif_canopy:units = "meters" ;
      	float h_max_canopy(delta_time) ;
      		h_max_canopy:_FillValue = 3.402823e+38f ;
      		h_max_canopy:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_max_canopy:description = "Relative maximum of individual canopy heights within segment. Relative canopy heights have been computed by differencing the canopy photon height from the estimated terrain surface. Should be equivalent to RH100 metric reported in the literature." ;
      		h_max_canopy:long_name = "maximum canopy height" ;
      		h_max_canopy:source = "Land ATBD section 2.2.12" ;
      		h_max_canopy:units = "meters" ;
      	float h_max_canopy_abs(delta_time) ;
      		h_max_canopy_abs:_FillValue = 3.402823e+38f ;
      		h_max_canopy_abs:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_max_canopy_abs:description = "Maximum of individual absolute canopy heights within segment referenced above the WGS84 ellipsoid." ;
      		h_max_canopy_abs:long_name = "absolute maximum canopy height" ;
      		h_max_canopy_abs:source = "Land ATBD section 2.2.11" ;
      		h_max_canopy_abs:units = "meters" ;
      	float h_mean_canopy(delta_time) ;
      		h_mean_canopy:_FillValue = 3.402823e+38f ;
      		h_mean_canopy:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_mean_canopy:description = "Mean of individual relative canopy heights within segment.  Relative canopy heights have been computed by differencing the canopy photon height from the estimated terrain surface." ;
      		h_mean_canopy:long_name = "mean canopy height" ;
      		h_mean_canopy:source = "Land ATBD section 4.12" ;
      		h_mean_canopy:units = "meters" ;
      	float h_mean_canopy_abs(delta_time) ;
      		h_mean_canopy_abs:_FillValue = 3.402823e+38f ;
      		h_mean_canopy_abs:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_mean_canopy_abs:description = "Mean of the individual absolute canopy heights within segment referenced above the WGS84 Ellipsoid." ;
      		h_mean_canopy_abs:long_name = "absolute mean canopy height" ;
      		h_mean_canopy_abs:source = "Land ATBD section 2.2.4" ;
      		h_mean_canopy_abs:units = "meters" ;
      	float h_median_canopy(delta_time) ;
      		h_median_canopy:_FillValue = 3.402823e+38f ;
      		h_median_canopy:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_median_canopy:description = "The median of individual relative canopy heights within segment. Relative canopy heights have been computed by differencing the canopy photon height from the estimated terrain surface. This parameter should be equivalent to RH50 reported in the literature." ;
      		h_median_canopy:long_name = "median canopy height" ;
      		h_median_canopy:source = "Land ATBD section 2.2.8" ;
      		h_median_canopy:units = "meters" ;
      	float h_median_canopy_abs(delta_time) ;
      		h_median_canopy_abs:_FillValue = 3.402823e+38f ;
      		h_median_canopy_abs:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_median_canopy_abs:description = "The median of individual absolute canopy heights within segment referenced above the WGS84 Ellipsoid." ;
      		h_median_canopy_abs:long_name = "absolute segment median canopy height" ;
      		h_median_canopy_abs:source = "Land ATBD section 2.2.6" ;
      		h_median_canopy_abs:units = "meters" ;
      	float h_min_canopy(delta_time) ;
      		h_min_canopy:_FillValue = 3.402823e+38f ;
      		h_min_canopy:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_min_canopy:description = "The minimum of relative individual canopy heights within segment. Relative canopy heights have been computed by differencing the canopy photon height from the estimated terrain surface." ;
      		h_min_canopy:long_name = "minimum canopy height" ;
      		h_min_canopy:source = "Land ATBD section 2.2.10" ;
      		h_min_canopy:units = "meters" ;
      	float h_min_canopy_abs(delta_time) ;
      		h_min_canopy_abs:_FillValue = 3.402823e+38f ;
      		h_min_canopy_abs:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_min_canopy_abs:description = "The minimum of absolute individual canopy heights within segment referenced above the WGS84 Ellipsoid." ;
      		h_min_canopy_abs:long_name = "absolute minimum canopy height" ;
      		h_min_canopy_abs:source = "Land ATBD section 2.2.9" ;
      		h_min_canopy_abs:units = "meters" ;
      	int landsat_flag(delta_time) ;
      		landsat_flag:_FillValue = 2147483647 ;
      		landsat_flag:coordinates = "../delta_time ../latitude ../longitude" ;
      		landsat_flag:description = "Flag indicating that more than 50% of the Landsat Continuous Cover product have values > 100 for the L-Km segment.  Canopy is assumed present along the L-km segment if landsat_flag is 1." ;
      		landsat_flag:flag_meanings = "canopy_not_assumed_present canopy_assumed_present" ;
      		landsat_flag:flag_values = 0, 1 ;
      		landsat_flag:long_name = "landsat flag" ;
      		landsat_flag:source = "Land ATBD section 2.2.25" ;
      		landsat_flag:units = "1" ;
      	float landsat_perc(delta_time) ;
      		landsat_perc:_FillValue = 3.402823e+38f ;
      		landsat_perc:coordinates = "../delta_time ../latitude ../longitude" ;
      		landsat_perc:description = "Average percentage value of the valid (value <= 100) Landsat Tree Cover Continuous Fields product for each 100 m segment" ;
      		landsat_perc:long_name = "landsat percentage canopy" ;
      		landsat_perc:source = "Land ATBD section 2.2.24" ;
      		landsat_perc:units = "1" ;
      	int n_ca_photons(delta_time) ;
      		n_ca_photons:coordinates = "../delta_time ../latitude ../longitude" ;
      		n_ca_photons:description = "The number of photons classified as canopy within the segment." ;
      		n_ca_photons:long_name = "number canopy photons" ;
      		n_ca_photons:source = "Land ATBD section 4.12" ;
      		n_ca_photons:units = "1" ;
      	int n_toc_photons(delta_time) ;
      		n_toc_photons:coordinates = "../delta_time ../latitude ../longitude" ;
      		n_toc_photons:description = "The number of photons classified as top of canopy within the segment." ;
      		n_toc_photons:long_name = "number top of canopy photons" ;
      		n_toc_photons:source = "Land ATBD section 4.12" ;
      		n_toc_photons:units = "1" ;
      	byte subset_can_flag(delta_time, ds_geosegments) ;
      		subset_can_flag:_FillValue = 127b ;
      		subset_can_flag:contentType = "modelResult" ;
      		subset_can_flag:coordinates = "../delta_time ../latitude ../longitude" ;
      		subset_can_flag:description = "Quality flag indicating the canopy photons populating the 100 m segment statistics are derived from less than 100 m worth of photons and/or less than 5 20m ATL03 segments." ;
      		subset_can_flag:flag_meanings = "no_photon_data_within_geosegment no_canopy_photons_within_geosegment canopy_photons_present_within_geosegment" ;
      		subset_can_flag:flag_values = -1b, 0b, 1b ;
      		subset_can_flag:long_name = "subset canopy flag" ;
      		subset_can_flag:source = "Land/Veg ATBD 15 Novemebr 2019, Section 2.2.25" ;
      		subset_can_flag:units = "1" ;
      		subset_can_flag:valid_max = 1b ;
      		subset_can_flag:valid_min = -1b ;
      	float toc_roughness(delta_time) ;
      		toc_roughness:_FillValue = 3.402823e+38f ;
      		toc_roughness:coordinates = "../delta_time ../latitude ../longitude" ;
      		toc_roughness:description = "Standard deviation of the relative heights of all photons classified as top of canopy within the segment" ;
      		toc_roughness:long_name = "top of canopy roughness" ;
      		toc_roughness:source = "Land ATBD section 4.12" ;
      		toc_roughness:units = "meters" ;

      // group attributes:
      		:Description = "Contains height parameters based on the land algorithm." ;
      		:data_rate = "Data are stored as aggregates of 100 meters." ;
      } // group canopy

    group: terrain {
      variables:
      	float h_te_best_fit(delta_time) ;
      		h_te_best_fit:_FillValue = 3.402823e+38f ;
      		h_te_best_fit:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_te_best_fit:description = "The best fit terrain elevation at the the mid-point location of each 100m segment. The mid-segment terrain elevation is determined by selecting the best of three fits- linear, 3rd order and 4th order polynomials - to the terrain photons and interpolating the elevation at the mid-point location of the 100 m segment. For the linear fit, a slope correction and weighting is applied to each ground photon based on the distance to the slope height at the center of the segment." ;
      		h_te_best_fit:long_name = "segment terrain height best fit" ;
      		h_te_best_fit:source = "Land ATBD section 2.1.15" ;
      		h_te_best_fit:units = "meters" ;
      	float h_te_interp(delta_time) ;
      		h_te_interp:_FillValue = 3.402823e+38f ;
      		h_te_interp:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_te_interp:description = "Interpolated terrain surface height above the WGS84 Ellipsoid at the midpoint of the segment." ;
      		h_te_interp:long_name = "interpolated terrain surface height" ;
      		h_te_interp:source = "Land ATBD section 4.9" ;
      		h_te_interp:units = "meters" ;
      	float h_te_max(delta_time) ;
      		h_te_max:_FillValue = 3.402823e+38f ;
      		h_te_max:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_te_max:description = "The maximum of the photon heights above the WGS84 Ellipsoid, classified as terrain within the segment." ;
      		h_te_max:long_name = "maximum terrain height" ;
      		h_te_max:source = "Land ATBD section 4.11" ;
      		h_te_max:units = "meters" ;
      	float h_te_mean(delta_time) ;
      		h_te_mean:_FillValue = 3.402823e+38f ;
      		h_te_mean:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_te_mean:description = "The mean of the photon heights above the WGS84 Ellipsoid, classified as terrain within the segment." ;
      		h_te_mean:long_name = "mean terrain height" ;
      		h_te_mean:source = "Land ATBD section 4.11" ;
      		h_te_mean:units = "meters" ;
      	float h_te_median(delta_time) ;
      		h_te_median:_FillValue = 3.402823e+38f ;
      		h_te_median:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_te_median:description = "The median of the photon heights above the WGS84 Ellipsoid, classified as terrain within the segment." ;
      		h_te_median:long_name = "median terrain height" ;
      		h_te_median:source = "Land ATBD section 4.11" ;
      		h_te_median:units = "meters" ;
      	float h_te_min(delta_time) ;
      		h_te_min:_FillValue = 3.402823e+38f ;
      		h_te_min:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_te_min:description = "The minimum of the photon heights above the WGS84 Ellipsoid, classified as terrain within the segment." ;
      		h_te_min:long_name = "minimum terrain height" ;
      		h_te_min:source = "Land ATBD section 4.11" ;
      		h_te_min:units = "meters" ;
      	float h_te_mode(delta_time) ;
      		h_te_mode:_FillValue = 3.402823e+38f ;
      		h_te_mode:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_te_mode:description = "The mode of the photon heights above the WGS84 Ellipsoid, classified as terrain within the segment." ;
      		h_te_mode:long_name = "mode of terrain heights" ;
      		h_te_mode:source = "Land ATBD section 4.11" ;
      		h_te_mode:units = "meters" ;
      	float h_te_skew(delta_time) ;
      		h_te_skew:_FillValue = 3.402823e+38f ;
      		h_te_skew:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_te_skew:description = "The skewness of the photon heights above the WGS84 Ellipsoid, classified as terrain within the segment." ;
      		h_te_skew:long_name = "skew of terrain heights" ;
      		h_te_skew:source = "Land ATBD section 4.11" ;
      		h_te_skew:units = "meters" ;
      	float h_te_std(delta_time) ;
      		h_te_std:_FillValue = 3.402823e+38f ;
      		h_te_std:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_te_std:description = "The standard deviation of the photon heights above the WGS84 Ellipsoid, classified as terrain within the segment." ;
      		h_te_std:long_name = "segment terrain roughness" ;
      		h_te_std:source = "Land ATBD section 4.11" ;
      		h_te_std:units = "meters" ;
      	float h_te_uncertainty(delta_time) ;
      		h_te_uncertainty:_FillValue = 3.402823e+38f ;
      		h_te_uncertainty:coordinates = "../delta_time ../latitude ../longitude" ;
      		h_te_uncertainty:description = "Uncertainty of the mean terrain height for the segment. This uncertainty incorporates all systematic uncertainties(e.g. timing orbits, geolocation,etc.) as well as uncertainty from errors of identified photons.  This parameter is described in section 1, equation 1.4" ;
      		h_te_uncertainty:long_name = "uncertainty of h_te_mean" ;
      		h_te_uncertainty:source = "Land ATBD section 4.11" ;
      		h_te_uncertainty:units = "meters" ;
      	int n_te_photons(delta_time) ;
      		n_te_photons:coordinates = "../delta_time ../latitude ../longitude" ;
      		n_te_photons:description = "The number of the photons classified as terrain within the segment." ;
      		n_te_photons:long_name = "number of ground photons" ;
      		n_te_photons:source = "Land ATBD section 4.11" ;
      		n_te_photons:units = "1" ;
      	byte subset_te_flag(delta_time, ds_geosegments) ;
      		subset_te_flag:_FillValue = 127b ;
      		subset_te_flag:contentType = "modelResult" ;
      		subset_te_flag:coordinates = "../delta_time ../latitude ../longitude" ;
      		subset_te_flag:description = "Quality flag indicating the terrain photons populating the 100 m segment statistics are derived from less than 100 m worth of photons and/or less than 5 20m ATL03 segments." ;
      		subset_te_flag:flag_meanings = "no_photon_data_within_geosegment no_terrain_photons_within_geosegment terrain_photons_present_within_geosegment" ;
      		subset_te_flag:flag_values = -1b, 0b, 1b ;
      		subset_te_flag:long_name = "subset terrain flag" ;
      		subset_te_flag:source = "Land/Veg ATBD 15 Novemebr 2019, Section 2.1.15" ;
      		subset_te_flag:units = "1" ;
      		subset_te_flag:valid_max = 1b ;
      		subset_te_flag:valid_min = -1b ;
      	float terrain_slope(delta_time) ;
      		terrain_slope:_FillValue = 3.402823e+38f ;
      		terrain_slope:coordinates = "../delta_time ../latitude ../longitude" ;
      		terrain_slope:description = "The along-track slope of terrain, within each segment;computed by a linear fit of terrain classified photons. Slope is in units of delta height over delta along track distance." ;
      		terrain_slope:long_name = "segment terrain slope" ;
      		terrain_slope:source = "Land ATBD section 4.11" ;
      		terrain_slope:units = "1" ;

      // group attributes:
      		:Description = "Contains terrain parameters at a 100m aggregation." ;
      		:data_rate = "Data are stored as aggregates of 100 meters." ;
      } // group terrain
    } // group land_segments
  } // group gt1r
}
